
module huffman_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module huffman_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_4 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_6 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman ( clk, reset, gray_valid, CNT_valid, gray_data, CNT1, CNT2, 
        CNT3, CNT4, CNT5, CNT6, code_valid, HC1, HC2, HC3, HC4, HC5, HC6, M1, 
        M2, M3, M4, M5, M6 );
  input [7:0] gray_data;
  output [7:0] CNT1;
  output [7:0] CNT2;
  output [7:0] CNT3;
  output [7:0] CNT4;
  output [7:0] CNT5;
  output [7:0] CNT6;
  output [7:0] HC1;
  output [7:0] HC2;
  output [7:0] HC3;
  output [7:0] HC4;
  output [7:0] HC5;
  output [7:0] HC6;
  output [7:0] M1;
  output [7:0] M2;
  output [7:0] M3;
  output [7:0] M4;
  output [7:0] M5;
  output [7:0] M6;
  input clk, reset, gray_valid;
  output CNT_valid, code_valid;
  wire   \SET[0][7] , \SET[0][6] , \SET[0][5] , \SET[0][4] , \SET[0][3] ,
         \SET[0][2] , \SET[0][1] , \SET[0][0] , \SET[1][7] , \SET[1][6] ,
         \SET[1][5] , \SET[1][4] , \SET[1][3] , \SET[1][2] , \SET[1][1] ,
         \SET[1][0] , \SET[2][7] , \SET[2][6] , \SET[2][5] , \SET[2][4] ,
         \SET[2][3] , \SET[2][2] , \SET[2][1] , \SET[2][0] , \SET[3][7] ,
         \SET[3][6] , \SET[3][5] , \SET[3][4] , \SET[3][3] , \SET[3][2] ,
         \SET[3][1] , \SET[3][0] , \SET[4][7] , \SET[4][6] , \SET[4][5] ,
         \SET[4][4] , \SET[4][3] , \SET[4][2] , \SET[4][1] , \SET[4][0] ,
         \SET[5][7] , \SET[5][6] , \SET[5][5] , \SET[5][4] , \SET[5][3] ,
         \SET[5][2] , \SET[5][1] , \SET[5][0] , N807, N808, N809, N810, N811,
         N812, N813, N814, N821, N822, N823, N824, N825, N826, N827, N828,
         \bitpos[0][2] , \bitpos[0][1] , \bitpos[0][0] , \bitpos[1][2] ,
         \bitpos[1][1] , \bitpos[1][0] , \bitpos[2][2] , \bitpos[2][1] ,
         \bitpos[2][0] , \bitpos[3][2] , \bitpos[3][1] , \bitpos[3][0] ,
         \bitpos[4][2] , \bitpos[4][1] , \bitpos[4][0] , \bitpos[5][2] ,
         \bitpos[5][1] , \bitpos[5][0] , \SET_flag[0][5] , \SET_flag[0][4] ,
         \SET_flag[0][3] , \SET_flag[0][2] , \SET_flag[0][1] ,
         \SET_flag[0][0] , \SET_flag[1][5] , \SET_flag[1][4] ,
         \SET_flag[1][3] , \SET_flag[1][2] , \SET_flag[1][1] ,
         \SET_flag[1][0] , \SET_flag[2][5] , \SET_flag[2][4] ,
         \SET_flag[2][3] , \SET_flag[2][2] , \SET_flag[2][1] ,
         \SET_flag[2][0] , \SET_flag[3][5] , \SET_flag[3][4] ,
         \SET_flag[3][3] , \SET_flag[3][2] , \SET_flag[3][1] ,
         \SET_flag[3][0] , \SET_flag[4][5] , \SET_flag[4][4] ,
         \SET_flag[4][3] , \SET_flag[4][2] , \SET_flag[4][1] ,
         \SET_flag[4][0] , \SET_flag[5][5] , \SET_flag[5][4] ,
         \SET_flag[5][3] , \SET_flag[5][2] , \SET_flag[5][1] ,
         \SET_flag[5][0] , N835, N836, N837, N838, N839, N840, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N947, N948, N949, N950, N951, N952, N953, N962, N1777,
         N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787,
         N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797,
         N1798, N1799, N1800, N1867, N1868, N1869, N1870, N1871, N1872, n68,
         n69, n81, n83, n84, n85, n86, n87, n88, n89, n90, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n472, n473,
         n474, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;
  wire   [2:0] state;
  wire   [2:0] nextstate;
  wire   [6:0] amount;
  wire   [2:0] times;
  wire   [2:0] endpoint;
  wire   [2:0] num;
  wire   [2:0] count;

  OAI211X2 U390 ( .A0(n1271), .A1(n405), .B0(n468), .C0(n469), .Y(n380) );
  OAI211X2 U397 ( .A0(n1277), .A1(n405), .B0(n478), .C0(n479), .Y(n385) );
  OAI211X2 U406 ( .A0(n1283), .A1(n405), .B0(n483), .C0(n484), .Y(n389) );
  OAI211X2 U415 ( .A0(n1289), .A1(n405), .B0(n488), .C0(n489), .Y(n393) );
  OAI211X2 U424 ( .A0(n1295), .A1(n405), .B0(n493), .C0(n494), .Y(n397) );
  OAI211X2 U437 ( .A0(n1301), .A1(n405), .B0(n500), .C0(n501), .Y(n406) );
  OAI221X2 U501 ( .A0(n541), .A1(n542), .B0(n192), .B1(n528), .C0(n1162), .Y(
        n425) );
  OAI211X2 U525 ( .A0(n556), .A1(n542), .B0(n1163), .C0(n557), .Y(n555) );
  OAI221X2 U553 ( .A0(n573), .A1(n542), .B0(n192), .B1(n559), .C0(n1162), .Y(
        n572) );
  OAI211X2 U579 ( .A0(n588), .A1(n542), .B0(n589), .C0(n1162), .Y(n587) );
  OAI211X2 U591 ( .A0(n192), .A1(n596), .B0(n1162), .C0(n597), .Y(n378) );
  OAI211X2 U718 ( .A0(n1266), .A1(n90), .B0(n645), .C0(n646), .Y(N828) );
  OAI211X2 U721 ( .A0(n1266), .A1(n89), .B0(n647), .C0(n648), .Y(N827) );
  OAI211X2 U724 ( .A0(n1266), .A1(n88), .B0(n649), .C0(n650), .Y(N826) );
  OAI211X2 U727 ( .A0(n1266), .A1(n87), .B0(n651), .C0(n652), .Y(N825) );
  OAI211X2 U730 ( .A0(n1266), .A1(n86), .B0(n653), .C0(n654), .Y(N824) );
  OAI211X2 U733 ( .A0(n1266), .A1(n85), .B0(n655), .C0(n656), .Y(N823) );
  OAI211X2 U739 ( .A0(n1266), .A1(n83), .B0(n659), .C0(n660), .Y(N821) );
  OAI211X2 U769 ( .A0(n405), .A1(n83), .B0(n675), .C0(n676), .Y(N807) );
  huffman_DW01_add_0 add_231 ( .A({N1777, N1778, N1779, N1780, N1781, N1782, 
        N1783, N1784}), .B({N1792, N1791, N1790, N1789, N1788, N1787, N1786, 
        N1785}), .CI(1'b0), .SUM({N1800, N1799, N1798, N1797, N1796, N1795, 
        N1794, N1793}) );
  huffman_DW01_inc_0 add_125 ( .A(amount), .SUM({N953, N952, N951, N950, N949, 
        N948, N947}) );
  huffman_DW01_inc_1 add_123 ( .A(CNT6), .SUM({N939, N938, N937, N936, N935, 
        N934, N933, N932}) );
  huffman_DW01_inc_2 add_122 ( .A(CNT5), .SUM({N931, N930, N929, N928, N927, 
        N926, N925, N924}) );
  huffman_DW01_inc_3 add_121 ( .A(CNT4), .SUM({N923, N922, N921, N920, N919, 
        N918, N917, N916}) );
  huffman_DW01_inc_4 add_120 ( .A(CNT3), .SUM({N915, N914, N913, N912, N911, 
        N910, N909, N908}) );
  huffman_DW01_inc_5 add_119 ( .A(CNT2), .SUM({N907, N906, N905, N904, N903, 
        N902, N901, N900}) );
  huffman_DW01_inc_6 add_118 ( .A(CNT1), .SUM({N899, N898, N897, N896, N895, 
        N894, N893, N892}) );
  DFFQX1 \amount_reg[6]  ( .D(n910), .CK(clk), .Q(amount[6]) );
  DFFQX1 \bitpos_reg[5][1]  ( .D(n789), .CK(clk), .Q(\bitpos[5][1] ) );
  DFFQX1 \bitpos_reg[4][1]  ( .D(n786), .CK(clk), .Q(\bitpos[4][1] ) );
  DFFQX1 \bitpos_reg[3][1]  ( .D(n783), .CK(clk), .Q(\bitpos[3][1] ) );
  DFFQX1 \bitpos_reg[2][1]  ( .D(n780), .CK(clk), .Q(\bitpos[2][1] ) );
  DFFQX1 \bitpos_reg[1][1]  ( .D(n777), .CK(clk), .Q(\bitpos[1][1] ) );
  DFFQX1 \bitpos_reg[0][1]  ( .D(n774), .CK(clk), .Q(\bitpos[0][1] ) );
  DFFQX1 \bitpos_reg[5][2]  ( .D(n788), .CK(clk), .Q(\bitpos[5][2] ) );
  DFFQX1 \bitpos_reg[4][2]  ( .D(n785), .CK(clk), .Q(\bitpos[4][2] ) );
  DFFQX1 \bitpos_reg[3][2]  ( .D(n782), .CK(clk), .Q(\bitpos[3][2] ) );
  DFFQX1 \bitpos_reg[2][2]  ( .D(n779), .CK(clk), .Q(\bitpos[2][2] ) );
  DFFQX1 \bitpos_reg[1][2]  ( .D(n776), .CK(clk), .Q(\bitpos[1][2] ) );
  DFFQX1 \bitpos_reg[0][2]  ( .D(n791), .CK(clk), .Q(\bitpos[0][2] ) );
  DFFQX1 \bitpos_reg[5][0]  ( .D(n790), .CK(clk), .Q(\bitpos[5][0] ) );
  DFFQX1 \bitpos_reg[4][0]  ( .D(n787), .CK(clk), .Q(\bitpos[4][0] ) );
  DFFQX1 \bitpos_reg[3][0]  ( .D(n784), .CK(clk), .Q(\bitpos[3][0] ) );
  DFFQX1 \bitpos_reg[2][0]  ( .D(n781), .CK(clk), .Q(\bitpos[2][0] ) );
  DFFQX1 \bitpos_reg[1][0]  ( .D(n778), .CK(clk), .Q(\bitpos[1][0] ) );
  DFFQX1 \bitpos_reg[0][0]  ( .D(n775), .CK(clk), .Q(\bitpos[0][0] ) );
  DFFQX1 \amount_reg[3]  ( .D(n906), .CK(clk), .Q(amount[3]) );
  DFFQX1 \amount_reg[4]  ( .D(n905), .CK(clk), .Q(amount[4]) );
  DFFQX1 \amount_reg[1]  ( .D(n908), .CK(clk), .Q(amount[1]) );
  DFFQX1 \amount_reg[5]  ( .D(n904), .CK(clk), .Q(amount[5]) );
  DFFQX1 \amount_reg[2]  ( .D(n907), .CK(clk), .Q(amount[2]) );
  DFFQX1 \amount_reg[0]  ( .D(n909), .CK(clk), .Q(amount[0]) );
  DFFQX2 \CNT2_reg[7]  ( .D(n863), .CK(clk), .Q(CNT2[7]) );
  DFFQX2 \CNT1_reg[7]  ( .D(n871), .CK(clk), .Q(CNT1[7]) );
  DFFQX1 \SET_flag_reg[0][5]  ( .D(n792), .CK(clk), .Q(\SET_flag[0][5] ) );
  DFFQX1 \SET_flag_reg[0][4]  ( .D(n793), .CK(clk), .Q(\SET_flag[0][4] ) );
  DFFQX1 \SET_flag_reg[0][3]  ( .D(n794), .CK(clk), .Q(\SET_flag[0][3] ) );
  DFFQX1 \SET_flag_reg[0][2]  ( .D(n795), .CK(clk), .Q(\SET_flag[0][2] ) );
  DFFQX1 \SET_flag_reg[0][1]  ( .D(n796), .CK(clk), .Q(\SET_flag[0][1] ) );
  DFFQX1 \SET_flag_reg[0][0]  ( .D(n797), .CK(clk), .Q(\SET_flag[0][0] ) );
  DFFQX1 \SET_flag_reg[2][5]  ( .D(n798), .CK(clk), .Q(\SET_flag[2][5] ) );
  DFFQX1 \SET_flag_reg[2][4]  ( .D(n799), .CK(clk), .Q(\SET_flag[2][4] ) );
  DFFQX1 \SET_flag_reg[2][3]  ( .D(n800), .CK(clk), .Q(\SET_flag[2][3] ) );
  DFFQX1 \SET_flag_reg[2][2]  ( .D(n801), .CK(clk), .Q(\SET_flag[2][2] ) );
  DFFQX1 \SET_flag_reg[2][1]  ( .D(n802), .CK(clk), .Q(\SET_flag[2][1] ) );
  DFFQX1 \SET_flag_reg[2][0]  ( .D(n803), .CK(clk), .Q(\SET_flag[2][0] ) );
  DFFQX1 \endpoint_reg[0]  ( .D(n912), .CK(clk), .Q(endpoint[0]) );
  DFFQX1 \endpoint_reg[2]  ( .D(n913), .CK(clk), .Q(endpoint[2]) );
  DFFQX1 \times_reg[1]  ( .D(n914), .CK(clk), .Q(times[1]) );
  DFFQX1 \times_reg[2]  ( .D(n916), .CK(clk), .Q(times[2]) );
  DFFX1 \SET_reg[0][6]  ( .D(n804), .CK(clk), .Q(\SET[0][6] ), .QN(n84) );
  DFFX1 \SET_reg[0][7]  ( .D(n852), .CK(clk), .Q(\SET[0][7] ), .QN(n83) );
  DFFQX1 \SET_reg[2][7]  ( .D(n819), .CK(clk), .Q(\SET[2][7] ) );
  DFFQX1 \SET_reg[4][7]  ( .D(n835), .CK(clk), .Q(\SET[4][7] ) );
  DFFQX1 \SET_reg[1][7]  ( .D(n811), .CK(clk), .Q(\SET[1][7] ) );
  DFFQX1 \SET_reg[5][7]  ( .D(n843), .CK(clk), .Q(\SET[5][7] ) );
  DFFX1 \SET_reg[0][0]  ( .D(n810), .CK(clk), .Q(\SET[0][0] ), .QN(n90) );
  DFFQX1 \SET_reg[2][0]  ( .D(n826), .CK(clk), .Q(\SET[2][0] ) );
  DFFQX1 \SET_reg[2][6]  ( .D(n820), .CK(clk), .Q(\SET[2][6] ) );
  DFFQX1 \SET_reg[4][6]  ( .D(n836), .CK(clk), .Q(\SET[4][6] ) );
  DFFQX1 \SET_reg[1][0]  ( .D(n818), .CK(clk), .Q(\SET[1][0] ) );
  DFFQX1 \SET_reg[1][3]  ( .D(n815), .CK(clk), .Q(\SET[1][3] ) );
  DFFQX1 \SET_reg[1][5]  ( .D(n813), .CK(clk), .Q(\SET[1][5] ) );
  DFFQX1 \SET_reg[1][6]  ( .D(n812), .CK(clk), .Q(\SET[1][6] ) );
  DFFQX1 \SET_reg[5][6]  ( .D(n844), .CK(clk), .Q(\SET[5][6] ) );
  DFFX1 \SET_reg[0][1]  ( .D(n809), .CK(clk), .Q(\SET[0][1] ), .QN(n89) );
  DFFX1 \SET_reg[0][2]  ( .D(n808), .CK(clk), .Q(\SET[0][2] ), .QN(n88) );
  DFFX1 \SET_reg[0][3]  ( .D(n807), .CK(clk), .Q(\SET[0][3] ), .QN(n87) );
  DFFX1 \SET_reg[0][4]  ( .D(n806), .CK(clk), .Q(\SET[0][4] ), .QN(n86) );
  DFFX1 \SET_reg[0][5]  ( .D(n805), .CK(clk), .Q(\SET[0][5] ), .QN(n85) );
  DFFQX1 \SET_reg[2][1]  ( .D(n825), .CK(clk), .Q(\SET[2][1] ) );
  DFFQX1 \SET_reg[2][2]  ( .D(n824), .CK(clk), .Q(\SET[2][2] ) );
  DFFQX1 \SET_reg[2][3]  ( .D(n823), .CK(clk), .Q(\SET[2][3] ) );
  DFFQX1 \SET_reg[2][4]  ( .D(n822), .CK(clk), .Q(\SET[2][4] ) );
  DFFQX1 \SET_reg[2][5]  ( .D(n821), .CK(clk), .Q(\SET[2][5] ) );
  DFFQX1 \SET_reg[4][0]  ( .D(n842), .CK(clk), .Q(\SET[4][0] ) );
  DFFQX1 \SET_reg[4][1]  ( .D(n841), .CK(clk), .Q(\SET[4][1] ) );
  DFFQX1 \SET_reg[4][2]  ( .D(n840), .CK(clk), .Q(\SET[4][2] ) );
  DFFQX1 \SET_reg[4][3]  ( .D(n839), .CK(clk), .Q(\SET[4][3] ) );
  DFFQX1 \SET_reg[4][4]  ( .D(n838), .CK(clk), .Q(\SET[4][4] ) );
  DFFQX1 \SET_reg[4][5]  ( .D(n837), .CK(clk), .Q(\SET[4][5] ) );
  DFFQX1 \SET_reg[1][1]  ( .D(n817), .CK(clk), .Q(\SET[1][1] ) );
  DFFQX1 \SET_reg[1][2]  ( .D(n816), .CK(clk), .Q(\SET[1][2] ) );
  DFFQX1 \SET_reg[1][4]  ( .D(n814), .CK(clk), .Q(\SET[1][4] ) );
  DFFQX1 \SET_reg[5][0]  ( .D(n850), .CK(clk), .Q(\SET[5][0] ) );
  DFFQX1 \SET_reg[5][1]  ( .D(n849), .CK(clk), .Q(\SET[5][1] ) );
  DFFQX1 \SET_reg[5][2]  ( .D(n848), .CK(clk), .Q(\SET[5][2] ) );
  DFFQX1 \SET_reg[5][3]  ( .D(n847), .CK(clk), .Q(\SET[5][3] ) );
  DFFQX1 \SET_reg[5][4]  ( .D(n846), .CK(clk), .Q(\SET[5][4] ) );
  DFFQX1 \SET_reg[5][5]  ( .D(n845), .CK(clk), .Q(\SET[5][5] ) );
  DFFQX2 \num_reg[0]  ( .D(n854), .CK(clk), .Q(num[0]) );
  DFFQX2 \CNT2_reg[2]  ( .D(n860), .CK(clk), .Q(CNT2[2]) );
  DFFQX2 \CNT2_reg[3]  ( .D(n859), .CK(clk), .Q(CNT2[3]) );
  DFFQX2 \CNT2_reg[4]  ( .D(n858), .CK(clk), .Q(CNT2[4]) );
  DFFQX2 \CNT2_reg[5]  ( .D(n857), .CK(clk), .Q(CNT2[5]) );
  DFFQX2 \CNT2_reg[6]  ( .D(n856), .CK(clk), .Q(CNT2[6]) );
  DFFQX2 \CNT1_reg[2]  ( .D(n868), .CK(clk), .Q(CNT1[2]) );
  DFFQX2 \CNT1_reg[3]  ( .D(n867), .CK(clk), .Q(CNT1[3]) );
  DFFQX2 \CNT1_reg[4]  ( .D(n866), .CK(clk), .Q(CNT1[4]) );
  DFFQX2 \CNT1_reg[5]  ( .D(n865), .CK(clk), .Q(CNT1[5]) );
  DFFQX2 \CNT1_reg[6]  ( .D(n864), .CK(clk), .Q(CNT1[6]) );
  DFFQX2 \CNT2_reg[1]  ( .D(n861), .CK(clk), .Q(CNT2[1]) );
  DFFQX2 \CNT1_reg[1]  ( .D(n869), .CK(clk), .Q(CNT1[1]) );
  DFFQX2 \CNT3_reg[1]  ( .D(n901), .CK(clk), .Q(CNT3[1]) );
  DFFQX2 \CNT2_reg[0]  ( .D(n862), .CK(clk), .Q(CNT2[0]) );
  DFFQX2 \CNT1_reg[0]  ( .D(n870), .CK(clk), .Q(CNT1[0]) );
  DFFQX2 \CNT3_reg[0]  ( .D(n902), .CK(clk), .Q(CNT3[0]) );
  DFFRX1 \state_reg[0]  ( .D(nextstate[0]), .CK(clk), .RN(n1162), .Q(state[0]), 
        .QN(n69) );
  DFFQX1 \times_reg[0]  ( .D(n915), .CK(clk), .Q(times[0]) );
  DFFRX1 \state_reg[1]  ( .D(nextstate[1]), .CK(clk), .RN(n1154), .Q(state[1])
         );
  DFFRX1 \state_reg[2]  ( .D(nextstate[2]), .CK(clk), .RN(n1162), .Q(state[2]), 
        .QN(n68) );
  DFFQX1 \SET_reg[3][7]  ( .D(n827), .CK(clk), .Q(\SET[3][7] ) );
  DFFQX1 \SET_reg[3][6]  ( .D(n828), .CK(clk), .Q(\SET[3][6] ) );
  DFFQX1 \SET_reg[3][0]  ( .D(n834), .CK(clk), .Q(\SET[3][0] ) );
  DFFQX1 \SET_reg[3][1]  ( .D(n833), .CK(clk), .Q(\SET[3][1] ) );
  DFFQX1 \SET_reg[3][2]  ( .D(n832), .CK(clk), .Q(\SET[3][2] ) );
  DFFQX1 \SET_reg[3][3]  ( .D(n831), .CK(clk), .Q(\SET[3][3] ) );
  DFFQX1 \SET_reg[3][4]  ( .D(n830), .CK(clk), .Q(\SET[3][4] ) );
  DFFQX1 \SET_reg[3][5]  ( .D(n829), .CK(clk), .Q(\SET[3][5] ) );
  EDFFTRX1 \endpoint_reg[1]  ( .RN(n1154), .D(n1261), .E(n1257), .CK(clk), .Q(
        endpoint[1]), .QN(n81) );
  DFFQX2 \num_reg[1]  ( .D(n851), .CK(clk), .Q(num[1]) );
  DFFQX2 \count_reg[0]  ( .D(n918), .CK(clk), .Q(count[0]) );
  DFFQX1 \count_reg[1]  ( .D(n855), .CK(clk), .Q(count[1]) );
  DFFQX1 \count_reg[2]  ( .D(n917), .CK(clk), .Q(count[2]) );
  EDFFX1 \SET_flag_reg[5][5]  ( .D(n1236), .E(n587), .CK(clk), .Q(
        \SET_flag[5][5] ) );
  EDFFX1 \SET_flag_reg[4][4]  ( .D(n1237), .E(n572), .CK(clk), .Q(
        \SET_flag[4][4] ) );
  EDFFX1 \SET_flag_reg[3][3]  ( .D(n1238), .E(n555), .CK(clk), .Q(
        \SET_flag[3][3] ) );
  EDFFX1 \SET_flag_reg[1][1]  ( .D(n1239), .E(n524), .CK(clk), .Q(
        \SET_flag[1][1] ), .QN(n1111) );
  EDFFX1 \SET_flag_reg[5][4]  ( .D(n1214), .E(n587), .CK(clk), .Q(
        \SET_flag[5][4] ) );
  EDFFX1 \SET_flag_reg[5][3]  ( .D(n1213), .E(n587), .CK(clk), .Q(
        \SET_flag[5][3] ) );
  EDFFX1 \SET_flag_reg[5][2]  ( .D(n1212), .E(n587), .CK(clk), .Q(
        \SET_flag[5][2] ) );
  EDFFX1 \SET_flag_reg[5][1]  ( .D(n1211), .E(n587), .CK(clk), .Q(
        \SET_flag[5][1] ) );
  EDFFX1 \SET_flag_reg[4][5]  ( .D(n1227), .E(n572), .CK(clk), .Q(
        \SET_flag[4][5] ) );
  EDFFX1 \SET_flag_reg[4][3]  ( .D(n1223), .E(n572), .CK(clk), .Q(
        \SET_flag[4][3] ) );
  EDFFX1 \SET_flag_reg[4][2]  ( .D(n1220), .E(n572), .CK(clk), .Q(
        \SET_flag[4][2] ) );
  EDFFX1 \SET_flag_reg[4][1]  ( .D(n1218), .E(n572), .CK(clk), .Q(
        \SET_flag[4][1] ) );
  EDFFX1 \SET_flag_reg[3][5]  ( .D(n1228), .E(n555), .CK(clk), .Q(
        \SET_flag[3][5] ) );
  EDFFX1 \SET_flag_reg[3][4]  ( .D(n1225), .E(n555), .CK(clk), .Q(
        \SET_flag[3][4] ) );
  EDFFX1 \SET_flag_reg[3][2]  ( .D(n1221), .E(n555), .CK(clk), .Q(
        \SET_flag[3][2] ) );
  EDFFX1 \SET_flag_reg[3][1]  ( .D(n1219), .E(n555), .CK(clk), .Q(
        \SET_flag[3][1] ) );
  EDFFX1 \SET_flag_reg[1][5]  ( .D(n1229), .E(n524), .CK(clk), .Q(
        \SET_flag[1][5] ), .QN(n1115) );
  EDFFX1 \SET_flag_reg[1][4]  ( .D(n1226), .E(n524), .CK(clk), .Q(
        \SET_flag[1][4] ), .QN(n1114) );
  EDFFX1 \SET_flag_reg[1][3]  ( .D(n1224), .E(n524), .CK(clk), .Q(
        \SET_flag[1][3] ), .QN(n1113) );
  EDFFX1 \SET_flag_reg[1][2]  ( .D(n1222), .E(n524), .CK(clk), .Q(
        \SET_flag[1][2] ), .QN(n1112) );
  EDFFX1 \SET_flag_reg[5][0]  ( .D(n1210), .E(n587), .CK(clk), .Q(
        \SET_flag[5][0] ) );
  EDFFX1 \SET_flag_reg[4][0]  ( .D(n1215), .E(n572), .CK(clk), .Q(
        \SET_flag[4][0] ) );
  EDFFX1 \SET_flag_reg[3][0]  ( .D(n1216), .E(n555), .CK(clk), .Q(
        \SET_flag[3][0] ) );
  EDFFX1 \SET_flag_reg[1][0]  ( .D(n1217), .E(n524), .CK(clk), .Q(
        \SET_flag[1][0] ), .QN(n1110) );
  DFFQX2 \CNT6_reg[0]  ( .D(n878), .CK(clk), .Q(CNT6[0]) );
  DFFQX2 \CNT5_reg[0]  ( .D(n886), .CK(clk), .Q(CNT5[0]) );
  DFFQX2 \CNT4_reg[0]  ( .D(n894), .CK(clk), .Q(CNT4[0]) );
  DFFQX2 \CNT6_reg[7]  ( .D(n879), .CK(clk), .Q(CNT6[7]) );
  DFFQX2 \CNT5_reg[7]  ( .D(n887), .CK(clk), .Q(CNT5[7]) );
  DFFQX2 \CNT4_reg[7]  ( .D(n895), .CK(clk), .Q(CNT4[7]) );
  DFFQX2 \CNT3_reg[7]  ( .D(n903), .CK(clk), .Q(CNT3[7]) );
  DFFQX2 \CNT6_reg[6]  ( .D(n872), .CK(clk), .Q(CNT6[6]) );
  DFFQX2 \CNT6_reg[5]  ( .D(n873), .CK(clk), .Q(CNT6[5]) );
  DFFQX2 \CNT6_reg[4]  ( .D(n874), .CK(clk), .Q(CNT6[4]) );
  DFFQX2 \CNT6_reg[3]  ( .D(n875), .CK(clk), .Q(CNT6[3]) );
  DFFQX2 \CNT6_reg[2]  ( .D(n876), .CK(clk), .Q(CNT6[2]) );
  DFFQX2 \CNT6_reg[1]  ( .D(n877), .CK(clk), .Q(CNT6[1]) );
  DFFQX2 \CNT5_reg[6]  ( .D(n880), .CK(clk), .Q(CNT5[6]) );
  DFFQX2 \CNT5_reg[5]  ( .D(n881), .CK(clk), .Q(CNT5[5]) );
  DFFQX2 \CNT5_reg[4]  ( .D(n882), .CK(clk), .Q(CNT5[4]) );
  DFFQX2 \CNT5_reg[3]  ( .D(n883), .CK(clk), .Q(CNT5[3]) );
  DFFQX2 \CNT5_reg[2]  ( .D(n884), .CK(clk), .Q(CNT5[2]) );
  DFFQX2 \CNT5_reg[1]  ( .D(n885), .CK(clk), .Q(CNT5[1]) );
  DFFQX2 \CNT4_reg[6]  ( .D(n888), .CK(clk), .Q(CNT4[6]) );
  DFFQX2 \CNT4_reg[5]  ( .D(n889), .CK(clk), .Q(CNT4[5]) );
  DFFQX2 \CNT4_reg[4]  ( .D(n890), .CK(clk), .Q(CNT4[4]) );
  DFFQX2 \CNT4_reg[3]  ( .D(n891), .CK(clk), .Q(CNT4[3]) );
  DFFQX2 \CNT4_reg[2]  ( .D(n892), .CK(clk), .Q(CNT4[2]) );
  DFFQX2 \CNT4_reg[1]  ( .D(n893), .CK(clk), .Q(CNT4[1]) );
  DFFQX2 \CNT3_reg[6]  ( .D(n896), .CK(clk), .Q(CNT3[6]) );
  DFFQX2 \CNT3_reg[5]  ( .D(n897), .CK(clk), .Q(CNT3[5]) );
  DFFQX2 \CNT3_reg[4]  ( .D(n898), .CK(clk), .Q(CNT3[4]) );
  DFFQX2 \CNT3_reg[3]  ( .D(n899), .CK(clk), .Q(CNT3[3]) );
  DFFQX2 \CNT3_reg[2]  ( .D(n900), .CK(clk), .Q(CNT3[2]) );
  DFFQX2 code_valid_reg ( .D(n677), .CK(clk), .Q(code_valid) );
  DFFQX2 \HC6_reg[3]  ( .D(n729), .CK(clk), .Q(HC6[3]) );
  DFFQX2 \HC6_reg[2]  ( .D(n728), .CK(clk), .Q(HC6[2]) );
  DFFQX2 \HC6_reg[1]  ( .D(n727), .CK(clk), .Q(HC6[1]) );
  DFFQX2 \HC6_reg[4]  ( .D(n730), .CK(clk), .Q(HC6[4]) );
  DFFQX2 \HC6_reg[0]  ( .D(n726), .CK(clk), .Q(HC6[0]) );
  DFFQX2 \HC3_reg[3]  ( .D(n753), .CK(clk), .Q(HC3[3]) );
  DFFQX2 \HC2_reg[3]  ( .D(n761), .CK(clk), .Q(HC2[3]) );
  DFFQX2 \HC1_reg[3]  ( .D(n769), .CK(clk), .Q(HC1[3]) );
  DFFQX2 \HC2_reg[2]  ( .D(n760), .CK(clk), .Q(HC2[2]) );
  DFFQX2 \HC1_reg[2]  ( .D(n768), .CK(clk), .Q(HC1[2]) );
  DFFQX2 \HC3_reg[7]  ( .D(n757), .CK(clk), .Q(HC3[7]) );
  DFFQX2 \HC3_reg[6]  ( .D(n756), .CK(clk), .Q(HC3[6]) );
  DFFQX2 \HC3_reg[4]  ( .D(n754), .CK(clk), .Q(HC3[4]) );
  DFFQX2 \HC2_reg[7]  ( .D(n765), .CK(clk), .Q(HC2[7]) );
  DFFQX2 \HC1_reg[7]  ( .D(n773), .CK(clk), .Q(HC1[7]) );
  DFFQX2 \HC1_reg[6]  ( .D(n772), .CK(clk), .Q(HC1[6]) );
  DFFQX2 \HC1_reg[4]  ( .D(n770), .CK(clk), .Q(HC1[4]) );
  DFFQX2 \HC1_reg[0]  ( .D(n766), .CK(clk), .Q(HC1[0]) );
  DFFQX2 \HC3_reg[2]  ( .D(n752), .CK(clk), .Q(HC3[2]) );
  DFFQX2 \HC3_reg[1]  ( .D(n751), .CK(clk), .Q(HC3[1]) );
  DFFQX2 \HC2_reg[1]  ( .D(n759), .CK(clk), .Q(HC2[1]) );
  DFFQX2 \HC1_reg[1]  ( .D(n767), .CK(clk), .Q(HC1[1]) );
  DFFQX2 \HC4_reg[7]  ( .D(n749), .CK(clk), .Q(HC4[7]) );
  DFFQX2 \HC4_reg[6]  ( .D(n748), .CK(clk), .Q(HC4[6]) );
  DFFQX2 \HC4_reg[5]  ( .D(n747), .CK(clk), .Q(HC4[5]) );
  DFFQX2 \HC4_reg[4]  ( .D(n746), .CK(clk), .Q(HC4[4]) );
  DFFQX2 \HC3_reg[5]  ( .D(n755), .CK(clk), .Q(HC3[5]) );
  DFFQX2 \HC3_reg[0]  ( .D(n750), .CK(clk), .Q(HC3[0]) );
  DFFQX2 \HC2_reg[6]  ( .D(n764), .CK(clk), .Q(HC2[6]) );
  DFFQX2 \HC2_reg[5]  ( .D(n763), .CK(clk), .Q(HC2[5]) );
  DFFQX2 \HC2_reg[4]  ( .D(n762), .CK(clk), .Q(HC2[4]) );
  DFFQX2 \HC2_reg[0]  ( .D(n758), .CK(clk), .Q(HC2[0]) );
  DFFQX2 \HC1_reg[5]  ( .D(n771), .CK(clk), .Q(HC1[5]) );
  DFFQX2 \HC5_reg[3]  ( .D(n737), .CK(clk), .Q(HC5[3]) );
  DFFQX2 \HC4_reg[3]  ( .D(n745), .CK(clk), .Q(HC4[3]) );
  DFFQX2 \HC5_reg[2]  ( .D(n736), .CK(clk), .Q(HC5[2]) );
  DFFQX2 \HC5_reg[1]  ( .D(n735), .CK(clk), .Q(HC5[1]) );
  DFFQX2 \HC4_reg[2]  ( .D(n744), .CK(clk), .Q(HC4[2]) );
  DFFQX2 \HC4_reg[1]  ( .D(n743), .CK(clk), .Q(HC4[1]) );
  DFFQX2 \HC6_reg[7]  ( .D(n733), .CK(clk), .Q(HC6[7]) );
  DFFQX2 \HC6_reg[6]  ( .D(n732), .CK(clk), .Q(HC6[6]) );
  DFFQX2 \HC6_reg[5]  ( .D(n731), .CK(clk), .Q(HC6[5]) );
  DFFQX2 \HC5_reg[7]  ( .D(n741), .CK(clk), .Q(HC5[7]) );
  DFFQX2 \HC5_reg[6]  ( .D(n740), .CK(clk), .Q(HC5[6]) );
  DFFQX2 \HC5_reg[5]  ( .D(n739), .CK(clk), .Q(HC5[5]) );
  DFFQX2 \HC5_reg[4]  ( .D(n738), .CK(clk), .Q(HC5[4]) );
  DFFQX2 \HC5_reg[0]  ( .D(n734), .CK(clk), .Q(HC5[0]) );
  DFFQX2 \HC4_reg[0]  ( .D(n742), .CK(clk), .Q(HC4[0]) );
  DFFQX2 CNT_valid_reg ( .D(n911), .CK(clk), .Q(CNT_valid) );
  DFFQX2 \M6_reg[3]  ( .D(n681), .CK(clk), .Q(M6[3]) );
  DFFQX2 \M6_reg[2]  ( .D(n680), .CK(clk), .Q(M6[2]) );
  DFFQX2 \M6_reg[1]  ( .D(n679), .CK(clk), .Q(M6[1]) );
  DFFQX2 \M6_reg[4]  ( .D(n682), .CK(clk), .Q(M6[4]) );
  DFFQX2 \M6_reg[0]  ( .D(n678), .CK(clk), .Q(M6[0]) );
  DFFQX2 \M3_reg[3]  ( .D(n705), .CK(clk), .Q(M3[3]) );
  DFFQX2 \M2_reg[3]  ( .D(n713), .CK(clk), .Q(M2[3]) );
  DFFQX2 \M1_reg[3]  ( .D(n721), .CK(clk), .Q(M1[3]) );
  DFFQX2 \M2_reg[2]  ( .D(n712), .CK(clk), .Q(M2[2]) );
  DFFQX2 \M1_reg[2]  ( .D(n720), .CK(clk), .Q(M1[2]) );
  DFFQX2 \M3_reg[7]  ( .D(n709), .CK(clk), .Q(M3[7]) );
  DFFQX2 \M3_reg[6]  ( .D(n708), .CK(clk), .Q(M3[6]) );
  DFFQX2 \M3_reg[4]  ( .D(n706), .CK(clk), .Q(M3[4]) );
  DFFQX2 \M2_reg[7]  ( .D(n717), .CK(clk), .Q(M2[7]) );
  DFFQX2 \M1_reg[7]  ( .D(n725), .CK(clk), .Q(M1[7]) );
  DFFQX2 \M1_reg[6]  ( .D(n724), .CK(clk), .Q(M1[6]) );
  DFFQX2 \M1_reg[4]  ( .D(n722), .CK(clk), .Q(M1[4]) );
  DFFQX2 \M1_reg[0]  ( .D(n718), .CK(clk), .Q(M1[0]) );
  DFFQX2 \M3_reg[2]  ( .D(n704), .CK(clk), .Q(M3[2]) );
  DFFQX2 \M3_reg[1]  ( .D(n703), .CK(clk), .Q(M3[1]) );
  DFFQX2 \M2_reg[1]  ( .D(n711), .CK(clk), .Q(M2[1]) );
  DFFQX2 \M1_reg[1]  ( .D(n719), .CK(clk), .Q(M1[1]) );
  DFFQX2 \M4_reg[7]  ( .D(n701), .CK(clk), .Q(M4[7]) );
  DFFQX2 \M4_reg[6]  ( .D(n700), .CK(clk), .Q(M4[6]) );
  DFFQX2 \M4_reg[5]  ( .D(n699), .CK(clk), .Q(M4[5]) );
  DFFQX2 \M4_reg[4]  ( .D(n698), .CK(clk), .Q(M4[4]) );
  DFFQX2 \M3_reg[5]  ( .D(n707), .CK(clk), .Q(M3[5]) );
  DFFQX2 \M3_reg[0]  ( .D(n702), .CK(clk), .Q(M3[0]) );
  DFFQX2 \M2_reg[6]  ( .D(n716), .CK(clk), .Q(M2[6]) );
  DFFQX2 \M2_reg[5]  ( .D(n715), .CK(clk), .Q(M2[5]) );
  DFFQX2 \M2_reg[4]  ( .D(n714), .CK(clk), .Q(M2[4]) );
  DFFQX2 \M2_reg[0]  ( .D(n710), .CK(clk), .Q(M2[0]) );
  DFFQX2 \M1_reg[5]  ( .D(n723), .CK(clk), .Q(M1[5]) );
  DFFQX2 \M5_reg[3]  ( .D(n689), .CK(clk), .Q(M5[3]) );
  DFFQX2 \M4_reg[3]  ( .D(n697), .CK(clk), .Q(M4[3]) );
  DFFQX2 \M5_reg[2]  ( .D(n688), .CK(clk), .Q(M5[2]) );
  DFFQX2 \M5_reg[1]  ( .D(n687), .CK(clk), .Q(M5[1]) );
  DFFQX2 \M4_reg[2]  ( .D(n696), .CK(clk), .Q(M4[2]) );
  DFFQX2 \M4_reg[1]  ( .D(n695), .CK(clk), .Q(M4[1]) );
  DFFQX2 \M6_reg[7]  ( .D(n685), .CK(clk), .Q(M6[7]) );
  DFFQX2 \M6_reg[6]  ( .D(n684), .CK(clk), .Q(M6[6]) );
  DFFQX2 \M6_reg[5]  ( .D(n683), .CK(clk), .Q(M6[5]) );
  DFFQX2 \M5_reg[7]  ( .D(n693), .CK(clk), .Q(M5[7]) );
  DFFQX2 \M5_reg[6]  ( .D(n692), .CK(clk), .Q(M5[6]) );
  DFFQX2 \M5_reg[5]  ( .D(n691), .CK(clk), .Q(M5[5]) );
  DFFQX2 \M5_reg[4]  ( .D(n690), .CK(clk), .Q(M5[4]) );
  DFFQX2 \M5_reg[0]  ( .D(n686), .CK(clk), .Q(M5[0]) );
  DFFQX2 \M4_reg[0]  ( .D(n694), .CK(clk), .Q(M4[0]) );
  DFFQX1 \num_reg[2]  ( .D(n853), .CK(clk), .Q(num[2]) );
  NOR2X4 U1060 ( .A(n193), .B(n1140), .Y(n1059) );
  CLKXOR2X4 U1061 ( .A(n1138), .B(n1067), .Y(n1060) );
  NOR2X4 U1062 ( .A(n1252), .B(count[0]), .Y(n1061) );
  NAND2X2 U1063 ( .A(num[1]), .B(n1265), .Y(n1062) );
  NOR2X4 U1064 ( .A(n1060), .B(n1261), .Y(n1063) );
  OAI221XL U1065 ( .A0(n1125), .A1(n1186), .B0(n1178), .B1(n1177), .C0(n1176), 
        .Y(n1179) );
  INVX3 U1066 ( .A(n425), .Y(n1195) );
  NAND2BX2 U1067 ( .AN(n572), .B(n1256), .Y(n560) );
  NAND2BX2 U1068 ( .AN(n555), .B(n1256), .Y(n543) );
  NAND2BX2 U1069 ( .AN(n587), .B(n1256), .Y(n575) );
  OAI21XL U1070 ( .A0(n1246), .A1(n1124), .B0(n1243), .Y(n526) );
  NAND2X2 U1071 ( .A(n1065), .B(n526), .Y(n524) );
  NOR2X4 U1072 ( .A(n1263), .B(count[0]), .Y(n1064) );
  NAND2BX2 U1073 ( .AN(n605), .B(N962), .Y(n542) );
  OAI22XL U1074 ( .A0(n1174), .A1(n1173), .B0(n1172), .B1(n1184), .Y(n1177) );
  OA21XL U1075 ( .A0(n192), .A1(n525), .B0(n1163), .Y(n1065) );
  CLKINVX1 U1076 ( .A(N827), .Y(n1185) );
  CLKINVX1 U1077 ( .A(N823), .Y(n1183) );
  INVX3 U1078 ( .A(n574), .Y(n1264) );
  CLKINVX1 U1079 ( .A(N825), .Y(n1184) );
  AOI222XL U1080 ( .A0(\SET[3][4] ), .A1(n1267), .B0(\SET[5][4] ), .B1(n1268), 
        .C0(\SET[4][4] ), .C1(n1264), .Y(n654) );
  INVX3 U1081 ( .A(count[2]), .Y(n1263) );
  INVX3 U1082 ( .A(count[1]), .Y(n1252) );
  CLKINVX1 U1083 ( .A(num[0]), .Y(n1265) );
  CLKINVX3 U1084 ( .A(n457), .Y(n1251) );
  CLKINVX3 U1085 ( .A(n434), .Y(n1245) );
  NAND2BX2 U1086 ( .AN(n524), .B(n1256), .Y(n512) );
  NOR2BXL U1087 ( .AN(N810), .B(N824), .Y(n1175) );
  NOR2X2 U1088 ( .A(n192), .B(n1140), .Y(n527) );
  NAND2BXL U1089 ( .AN(N812), .B(N826), .Y(n1172) );
  NAND2XL U1090 ( .A(n1061), .B(n1263), .Y(n434) );
  NAND2XL U1091 ( .A(n1064), .B(n1252), .Y(n457) );
  OA21XL U1092 ( .A0(N840), .A1(n1126), .B0(n1257), .Y(n333) );
  OA21XL U1093 ( .A0(N839), .A1(n1131), .B0(n1257), .Y(n318) );
  OA21XL U1094 ( .A0(N838), .A1(n1130), .B0(n1257), .Y(n303) );
  OA21XL U1095 ( .A0(N837), .A1(n1129), .B0(n1257), .Y(n288) );
  OA21XL U1096 ( .A0(N836), .A1(n1128), .B0(n1257), .Y(n273) );
  OA21XL U1097 ( .A0(N835), .A1(n1127), .B0(n1257), .Y(n258) );
  NOR2X1 U1098 ( .A(n630), .B(n1257), .Y(n604) );
  CLKINVX1 U1099 ( .A(n403), .Y(n1259) );
  INVX1 U1100 ( .A(count[0]), .Y(n1244) );
  AOI2BB2XL U1101 ( .B0(\SET[2][7] ), .B1(n1061), .A0N(n420), .A1N(n1341), .Y(
        n675) );
  AOI2BB2XL U1102 ( .B0(\SET[2][6] ), .B1(n1061), .A0N(n420), .A1N(n1337), .Y(
        n673) );
  AOI2BB1XL U1103 ( .A0N(num[1]), .A1N(n574), .B0(n1251), .Y(n573) );
  AOI2BB1XL U1104 ( .A0N(num[2]), .A1N(n558), .B0(n1247), .Y(n556) );
  AOI2BB1XL U1105 ( .A0N(num[1]), .A1N(n590), .B0(n1249), .Y(n588) );
  AOI2BB2XL U1106 ( .B0(n1124), .B1(\SET[1][7] ), .A0N(n1342), .A1N(n1062), 
        .Y(n659) );
  NOR3XL U1107 ( .A(num[1]), .B(num[2]), .C(n1265), .Y(n474) );
  AOI2BB2XL U1108 ( .B0(n1253), .B1(n1208), .A0N(count[0]), .A1N(n601), .Y(
        n644) );
  NOR3X1 U1109 ( .A(num[1]), .B(num[2]), .C(num[0]), .Y(n598) );
  NAND3X2 U1110 ( .A(n1252), .B(n1263), .C(count[0]), .Y(n420) );
  AOI2BB2XL U1111 ( .B0(n1124), .B1(\SET[1][6] ), .A0N(n1338), .A1N(n1062), 
        .Y(n657) );
  NAND2XL U1112 ( .A(count[2]), .B(count[0]), .Y(n643) );
  NAND2XL U1113 ( .A(count[1]), .B(count[0]), .Y(n610) );
  AO22XL U1114 ( .A0(num[0]), .A1(n1205), .B0(n591), .B1(n603), .Y(n854) );
  XNOR2X1 U1115 ( .A(n81), .B(n1132), .Y(n377) );
  NAND3X1 U1116 ( .A(n69), .B(n68), .C(state[1]), .Y(n193) );
  AOI22XL U1117 ( .A0(n1061), .A1(\SET_flag[2][0] ), .B0(\SET_flag[1][0] ), 
        .B1(n1246), .Y(n500) );
  AOI22XL U1118 ( .A0(n1061), .A1(\SET_flag[2][1] ), .B0(\SET_flag[1][1] ), 
        .B1(n1246), .Y(n493) );
  AOI22XL U1119 ( .A0(n1061), .A1(\SET_flag[2][2] ), .B0(\SET_flag[1][2] ), 
        .B1(n1246), .Y(n488) );
  AOI22XL U1120 ( .A0(n1061), .A1(\SET_flag[2][3] ), .B0(\SET_flag[1][3] ), 
        .B1(n1246), .Y(n483) );
  AOI22XL U1121 ( .A0(n1061), .A1(\SET_flag[2][4] ), .B0(\SET_flag[1][4] ), 
        .B1(n1246), .Y(n478) );
  AOI22XL U1122 ( .A0(n1061), .A1(\SET_flag[2][5] ), .B0(\SET_flag[1][5] ), 
        .B1(n1246), .Y(n468) );
  AOI2BB2XL U1123 ( .B0(\SET_flag[1][1] ), .B1(n1124), .A0N(n1062), .A1N(n1294), .Y(n495) );
  AOI2BB2XL U1124 ( .B0(\SET_flag[1][2] ), .B1(n1124), .A0N(n1062), .A1N(n1288), .Y(n490) );
  AOI2BB2XL U1125 ( .B0(\SET_flag[1][3] ), .B1(n1124), .A0N(n1062), .A1N(n1282), .Y(n485) );
  AOI2BB2XL U1126 ( .B0(\SET_flag[1][4] ), .B1(n1124), .A0N(n1062), .A1N(n1276), .Y(n480) );
  AOI2BB2XL U1127 ( .B0(\SET_flag[1][5] ), .B1(n1124), .A0N(n1062), .A1N(n1270), .Y(n472) );
  OR2X1 U1128 ( .A(N1868), .B(N839), .Y(n398) );
  OR2X1 U1129 ( .A(N1869), .B(N838), .Y(n394) );
  OR2X1 U1130 ( .A(N1870), .B(N837), .Y(n390) );
  OR2X1 U1131 ( .A(N1871), .B(N836), .Y(n386) );
  OR2X1 U1132 ( .A(N1872), .B(N835), .Y(n382) );
  AOI2BB2XL U1133 ( .B0(\SET_flag[1][0] ), .B1(n1124), .A0N(n1062), .A1N(n1300), .Y(n498) );
  INVXL U1134 ( .A(num[1]), .Y(n1269) );
  NAND3X2 U1135 ( .A(state[0]), .B(n68), .C(state[1]), .Y(n192) );
  OAI211X4 U1136 ( .A0(n405), .A1(n86), .B0(n669), .C0(n670), .Y(N810) );
  OAI211X4 U1137 ( .A0(n405), .A1(n88), .B0(n665), .C0(n666), .Y(N812) );
  OAI211X4 U1138 ( .A0(n405), .A1(n89), .B0(n663), .C0(n664), .Y(N813) );
  OAI211X4 U1139 ( .A0(n405), .A1(n90), .B0(n661), .C0(n662), .Y(N814) );
  OAI211X4 U1140 ( .A0(n405), .A1(n84), .B0(n673), .C0(n674), .Y(N808) );
  INVX3 U1141 ( .A(n1066), .Y(n405) );
  INVX3 U1142 ( .A(n594), .Y(n1208) );
  CLKBUFX3 U1143 ( .A(n505), .Y(n1136) );
  CLKBUFX3 U1144 ( .A(n505), .Y(n1135) );
  CLKBUFX3 U1145 ( .A(n505), .Y(n1134) );
  NOR2BX2 U1146 ( .AN(n540), .B(n1245), .Y(n531) );
  AND2X2 U1147 ( .A(n1059), .B(n529), .Y(n540) );
  NOR2BX2 U1148 ( .AN(n571), .B(n1251), .Y(n562) );
  NOR2BX2 U1149 ( .AN(n554), .B(n1247), .Y(n545) );
  NOR2BX2 U1150 ( .AN(n586), .B(n1249), .Y(n577) );
  NAND2X1 U1151 ( .A(n1066), .B(n1059), .Y(n594) );
  INVX3 U1152 ( .A(n504), .Y(n1196) );
  INVX3 U1153 ( .A(n601), .Y(n1209) );
  INVX3 U1154 ( .A(n1161), .Y(n1140) );
  AND2XL U1155 ( .A(n1059), .B(n512), .Y(n523) );
  NOR2BX1 U1156 ( .AN(n1059), .B(n1249), .Y(n477) );
  NOR2BX1 U1157 ( .AN(n1059), .B(n1251), .Y(n452) );
  NOR2BX1 U1158 ( .AN(n1059), .B(n1247), .Y(n440) );
  NOR2BX1 U1159 ( .AN(n1059), .B(n1245), .Y(n427) );
  NAND2X1 U1160 ( .A(n1059), .B(n636), .Y(n635) );
  CLKINVX1 U1161 ( .A(n636), .Y(n1206) );
  NAND2X1 U1162 ( .A(n340), .B(n1160), .Y(n339) );
  NAND2X1 U1163 ( .A(n344), .B(n1154), .Y(n341) );
  NAND2X1 U1164 ( .A(n352), .B(n1159), .Y(n349) );
  NAND2X1 U1165 ( .A(n358), .B(n1158), .Y(n355) );
  NAND2X1 U1166 ( .A(n364), .B(n1161), .Y(n361) );
  NAND2X1 U1167 ( .A(n370), .B(n1159), .Y(n367) );
  CLKINVX1 U1168 ( .A(n462), .Y(n1232) );
  CLKINVX1 U1169 ( .A(n450), .Y(n1233) );
  CLKINVX1 U1170 ( .A(n424), .Y(n1235) );
  CLKINVX1 U1171 ( .A(n438), .Y(n1234) );
  CLKINVX1 U1172 ( .A(n606), .Y(n1207) );
  CLKINVX1 U1173 ( .A(n591), .Y(n1205) );
  INVX3 U1174 ( .A(n1158), .Y(n1143) );
  INVX3 U1175 ( .A(n1157), .Y(n1144) );
  INVX3 U1176 ( .A(n1156), .Y(n1145) );
  INVX3 U1177 ( .A(n1152), .Y(n1149) );
  INVX3 U1178 ( .A(n1155), .Y(n1146) );
  INVX3 U1179 ( .A(n1151), .Y(n1150) );
  INVX3 U1180 ( .A(n1154), .Y(n1147) );
  INVX3 U1181 ( .A(n1153), .Y(n1148) );
  INVX3 U1182 ( .A(n1160), .Y(n1141) );
  INVX3 U1183 ( .A(n1159), .Y(n1142) );
  CLKBUFX3 U1184 ( .A(n1132), .Y(n1121) );
  CLKBUFX3 U1185 ( .A(n1117), .Y(n1116) );
  NOR2BX2 U1186 ( .AN(n540), .B(n434), .Y(n532) );
  NAND2X2 U1187 ( .A(n1195), .B(n1256), .Y(n529) );
  CLKBUFX3 U1188 ( .A(n1164), .Y(n1162) );
  NOR2BX2 U1189 ( .AN(n523), .B(n1246), .Y(n514) );
  NOR2BX2 U1190 ( .AN(n571), .B(n457), .Y(n563) );
  NOR2BX2 U1191 ( .AN(n554), .B(n446), .Y(n546) );
  NOR2BX2 U1192 ( .AN(n586), .B(n467), .Y(n578) );
  NAND2X1 U1193 ( .A(n1059), .B(n405), .Y(n601) );
  NOR2X2 U1194 ( .A(n1203), .B(n1140), .Y(n624) );
  INVX3 U1195 ( .A(n381), .Y(n1230) );
  NAND2X2 U1196 ( .A(n1197), .B(n1256), .Y(n504) );
  CLKINVX1 U1197 ( .A(n542), .Y(n1243) );
  CLKBUFX3 U1198 ( .A(n1165), .Y(n1161) );
  CLKBUFX3 U1199 ( .A(n1164), .Y(n1163) );
  AND2XL U1200 ( .A(n1059), .B(n560), .Y(n571) );
  AND2XL U1201 ( .A(n1059), .B(n543), .Y(n554) );
  AND2XL U1202 ( .A(n1059), .B(n575), .Y(n586) );
  OAI211X1 U1203 ( .A0(n605), .A1(n405), .B0(n1163), .C0(n604), .Y(n636) );
  NOR2BX1 U1204 ( .AN(n1059), .B(n1246), .Y(n409) );
  AOI2BB1X1 U1205 ( .A0N(n251), .A1N(n252), .B0(n1143), .Y(n201) );
  AOI2BB1X1 U1206 ( .A0N(n266), .A1N(n267), .B0(n1144), .Y(n209) );
  AOI2BB1X1 U1207 ( .A0N(n281), .A1N(n282), .B0(n1144), .Y(n217) );
  AOI2BB1X1 U1208 ( .A0N(n296), .A1N(n297), .B0(n1145), .Y(n225) );
  AOI2BB1X1 U1209 ( .A0N(n311), .A1N(n312), .B0(n1145), .Y(n233) );
  AOI2BB1X1 U1210 ( .A0N(n326), .A1N(n327), .B0(n1146), .Y(n241) );
  AOI2BB1X1 U1211 ( .A0N(n252), .A1N(n1272), .B0(n1143), .Y(n204) );
  AOI2BB1X1 U1212 ( .A0N(n267), .A1N(n1278), .B0(n1144), .Y(n212) );
  AOI2BB1X1 U1213 ( .A0N(n282), .A1N(n1284), .B0(n1144), .Y(n220) );
  AOI2BB1X1 U1214 ( .A0N(n297), .A1N(n1290), .B0(n1146), .Y(n228) );
  AOI2BB1X1 U1215 ( .A0N(n312), .A1N(n1296), .B0(n1146), .Y(n236) );
  AOI2BB1X1 U1216 ( .A0N(n327), .A1N(n1302), .B0(n1146), .Y(n244) );
  NOR2X2 U1217 ( .A(n627), .B(n1140), .Y(n628) );
  NOR2X1 U1218 ( .A(n1256), .B(n1140), .Y(n505) );
  NAND2X1 U1219 ( .A(n1206), .B(n542), .Y(n591) );
  NAND2X2 U1220 ( .A(n456), .B(n527), .Y(n462) );
  NAND2X2 U1221 ( .A(n445), .B(n527), .Y(n450) );
  NAND2X2 U1222 ( .A(n419), .B(n527), .Y(n424) );
  NAND2X2 U1223 ( .A(n433), .B(n527), .Y(n438) );
  NAND2BX1 U1224 ( .AN(n333), .B(n1153), .Y(n340) );
  NAND2BX1 U1225 ( .AN(n318), .B(n1151), .Y(n344) );
  NAND2BX1 U1226 ( .AN(n303), .B(n1152), .Y(n352) );
  NAND2BX1 U1227 ( .AN(n288), .B(n1154), .Y(n358) );
  NAND2BX1 U1228 ( .AN(n273), .B(n1155), .Y(n364) );
  NAND2BX1 U1229 ( .AN(n258), .B(n1156), .Y(n370) );
  NAND3X1 U1230 ( .A(n605), .B(n1153), .C(n604), .Y(n606) );
  CLKINVX1 U1231 ( .A(n502), .Y(n1231) );
  OAI22XL U1232 ( .A0(n1133), .A1(n631), .B0(n1204), .B1(n632), .Y(n912) );
  NOR2X1 U1233 ( .A(n1140), .B(n1133), .Y(n632) );
  CLKINVX1 U1234 ( .A(n631), .Y(n1204) );
  CLKBUFX3 U1235 ( .A(n1167), .Y(n1153) );
  CLKBUFX3 U1236 ( .A(n1167), .Y(n1152) );
  CLKBUFX3 U1237 ( .A(n1167), .Y(n1154) );
  CLKBUFX3 U1238 ( .A(n1166), .Y(n1155) );
  CLKBUFX3 U1239 ( .A(n1167), .Y(n1151) );
  CLKBUFX3 U1240 ( .A(n1166), .Y(n1156) );
  CLKBUFX3 U1241 ( .A(n1166), .Y(n1157) );
  CLKBUFX3 U1242 ( .A(n1166), .Y(n1158) );
  CLKBUFX3 U1243 ( .A(n1165), .Y(n1160) );
  CLKBUFX3 U1244 ( .A(n1165), .Y(n1159) );
  NOR2X1 U1245 ( .A(n528), .B(n1133), .Y(n433) );
  INVX3 U1246 ( .A(n446), .Y(n1247) );
  INVX3 U1247 ( .A(n467), .Y(n1249) );
  CLKBUFX3 U1248 ( .A(endpoint[1]), .Y(n1119) );
  CLKBUFX3 U1249 ( .A(n1137), .Y(n1117) );
  CLKINVX1 U1250 ( .A(N1794), .Y(n1193) );
  CLKINVX1 U1251 ( .A(n369), .Y(n1272) );
  CLKINVX1 U1252 ( .A(n363), .Y(n1278) );
  CLKINVX1 U1253 ( .A(n357), .Y(n1284) );
  CLKINVX1 U1254 ( .A(n351), .Y(n1290) );
  CLKINVX1 U1255 ( .A(n343), .Y(n1296) );
  CLKINVX1 U1256 ( .A(n374), .Y(n1302) );
  CLKINVX1 U1257 ( .A(N821), .Y(n1182) );
  INVX3 U1258 ( .A(n610), .Y(n1248) );
  INVX3 U1259 ( .A(n643), .Y(n1250) );
  INVX3 U1260 ( .A(n598), .Y(n1266) );
  CLKINVX1 U1261 ( .A(n1139), .Y(n1164) );
  NAND2X1 U1262 ( .A(n377), .B(n1138), .Y(n525) );
  NOR2BX2 U1263 ( .AN(n523), .B(n420), .Y(n515) );
  INVX3 U1264 ( .A(n378), .Y(n1197) );
  NOR2BX2 U1265 ( .AN(n527), .B(n191), .Y(n381) );
  NOR2X2 U1266 ( .A(n1199), .B(n1140), .Y(n614) );
  NOR2X2 U1267 ( .A(n1198), .B(n1140), .Y(n611) );
  NOR2X2 U1268 ( .A(n1202), .B(n1140), .Y(n621) );
  NOR2X2 U1269 ( .A(n1201), .B(n1140), .Y(n619) );
  NOR2X2 U1270 ( .A(n1200), .B(n1140), .Y(n616) );
  INVX3 U1271 ( .A(n625), .Y(n1203) );
  OAI31XL U1272 ( .A0(n1242), .A1(n613), .A2(n1241), .B0(n1159), .Y(n625) );
  OAI22XL U1273 ( .A0(n1300), .A1(n425), .B0(n1195), .B1(n437), .Y(n803) );
  AOI222XL U1274 ( .A0(n1234), .A1(n1259), .B0(n427), .B1(n406), .C0(n1245), 
        .C1(n422), .Y(n437) );
  OAI22XL U1275 ( .A0(n1294), .A1(n425), .B0(n1195), .B1(n435), .Y(n802) );
  AOI222XL U1276 ( .A0(n1234), .A1(n398), .B0(n436), .B1(n1245), .C0(n427), 
        .C1(n397), .Y(n435) );
  OAI22XL U1277 ( .A0(n1288), .A1(n425), .B0(n1195), .B1(n430), .Y(n801) );
  AOI211X1 U1278 ( .A0(n1255), .A1(n431), .B0(n1149), .C0(n432), .Y(n430) );
  AND3X2 U1279 ( .A(n433), .B(n394), .C(n1257), .Y(n432) );
  AO22X1 U1280 ( .A0(n395), .A1(n1245), .B0(n434), .B1(n393), .Y(n431) );
  OAI22XL U1281 ( .A0(n1282), .A1(n425), .B0(n1195), .B1(n429), .Y(n800) );
  AOI222XL U1282 ( .A0(n1234), .A1(n390), .B0(n1245), .B1(n413), .C0(n427), 
        .C1(n389), .Y(n429) );
  OAI22XL U1283 ( .A0(n1276), .A1(n425), .B0(n1195), .B1(n428), .Y(n799) );
  AOI222XL U1284 ( .A0(n1234), .A1(n386), .B0(n1245), .B1(n411), .C0(n427), 
        .C1(n385), .Y(n428) );
  OAI22XL U1285 ( .A0(n1270), .A1(n425), .B0(n1195), .B1(n426), .Y(n798) );
  AOI222XL U1286 ( .A0(n1234), .A1(n382), .B0(n1245), .B1(n408), .C0(n427), 
        .C1(n380), .Y(n426) );
  OAI22XL U1287 ( .A0(n1301), .A1(n378), .B0(n1197), .B1(n400), .Y(n797) );
  AOI211X1 U1288 ( .A0(n1255), .A1(n401), .B0(n1149), .C0(n402), .Y(n400) );
  NOR3X1 U1289 ( .A(n192), .B(n403), .C(n191), .Y(n402) );
  AO22X1 U1290 ( .A0(n404), .A1(n1066), .B0(n405), .B1(n406), .Y(n401) );
  OAI22XL U1291 ( .A0(n1295), .A1(n378), .B0(n1197), .B1(n396), .Y(n796) );
  AOI222XL U1292 ( .A0(n1209), .A1(n397), .B0(n381), .B1(n398), .C0(n1208), 
        .C1(n399), .Y(n396) );
  OAI22XL U1293 ( .A0(n1289), .A1(n378), .B0(n1197), .B1(n392), .Y(n795) );
  AOI222XL U1294 ( .A0(n1209), .A1(n393), .B0(n381), .B1(n394), .C0(n1208), 
        .C1(n395), .Y(n392) );
  OAI22XL U1295 ( .A0(n1283), .A1(n378), .B0(n1197), .B1(n388), .Y(n794) );
  AOI222XL U1296 ( .A0(n1209), .A1(n389), .B0(n381), .B1(n390), .C0(n1208), 
        .C1(n391), .Y(n388) );
  OAI22XL U1297 ( .A0(n1277), .A1(n378), .B0(n1197), .B1(n384), .Y(n793) );
  AOI222XL U1298 ( .A0(n1209), .A1(n385), .B0(n381), .B1(n386), .C0(n1208), 
        .C1(n387), .Y(n384) );
  OAI22XL U1299 ( .A0(n1271), .A1(n378), .B0(n1197), .B1(n379), .Y(n792) );
  AOI222XL U1300 ( .A0(n1209), .A1(n380), .B0(n381), .B1(n382), .C0(n1208), 
        .C1(n383), .Y(n379) );
  INVX3 U1301 ( .A(n590), .Y(n1268) );
  INVX3 U1302 ( .A(n558), .Y(n1267) );
  AND3X2 U1303 ( .A(n1252), .B(n1263), .C(n1244), .Y(n1066) );
  CLKINVX1 U1304 ( .A(n1139), .Y(n1165) );
  CLKINVX1 U1305 ( .A(n461), .Y(n1215) );
  AOI222XL U1306 ( .A0(n1232), .A1(n1259), .B0(n452), .B1(n406), .C0(n1251), 
        .C1(n422), .Y(n461) );
  CLKINVX1 U1307 ( .A(n449), .Y(n1216) );
  AOI222XL U1308 ( .A0(n1233), .A1(n1259), .B0(n440), .B1(n406), .C0(n1247), 
        .C1(n422), .Y(n449) );
  CLKINVX1 U1309 ( .A(n421), .Y(n1217) );
  AOI222XL U1310 ( .A0(n1235), .A1(n1259), .B0(n409), .B1(n406), .C0(n422), 
        .C1(n1246), .Y(n421) );
  CLKINVX1 U1311 ( .A(n497), .Y(n1210) );
  AOI222XL U1312 ( .A0(n1231), .A1(n1259), .B0(n477), .B1(n406), .C0(n1249), 
        .C1(n422), .Y(n497) );
  CLKINVX1 U1313 ( .A(n460), .Y(n1218) );
  AOI222XL U1314 ( .A0(n1232), .A1(n398), .B0(n1251), .B1(n436), .C0(n452), 
        .C1(n397), .Y(n460) );
  CLKINVX1 U1315 ( .A(n448), .Y(n1219) );
  AOI222XL U1316 ( .A0(n1233), .A1(n398), .B0(n1247), .B1(n436), .C0(n440), 
        .C1(n397), .Y(n448) );
  CLKINVX1 U1317 ( .A(n492), .Y(n1211) );
  AOI222XL U1318 ( .A0(n1231), .A1(n398), .B0(n1249), .B1(n436), .C0(n477), 
        .C1(n397), .Y(n492) );
  CLKINVX1 U1319 ( .A(n459), .Y(n1220) );
  AOI222XL U1320 ( .A0(n1232), .A1(n394), .B0(n1251), .B1(n415), .C0(n452), 
        .C1(n393), .Y(n459) );
  CLKINVX1 U1321 ( .A(n447), .Y(n1221) );
  AOI222XL U1322 ( .A0(n1233), .A1(n394), .B0(n1247), .B1(n415), .C0(n440), 
        .C1(n393), .Y(n447) );
  CLKINVX1 U1323 ( .A(n487), .Y(n1212) );
  AOI222XL U1324 ( .A0(n1231), .A1(n394), .B0(n1249), .B1(n415), .C0(n477), 
        .C1(n393), .Y(n487) );
  CLKINVX1 U1325 ( .A(n458), .Y(n1223) );
  AOI222XL U1326 ( .A0(n1232), .A1(n390), .B0(n1251), .B1(n413), .C0(n452), 
        .C1(n389), .Y(n458) );
  CLKINVX1 U1327 ( .A(n482), .Y(n1213) );
  AOI222XL U1328 ( .A0(n1231), .A1(n390), .B0(n1249), .B1(n413), .C0(n477), 
        .C1(n389), .Y(n482) );
  CLKINVX1 U1329 ( .A(n441), .Y(n1225) );
  AOI222XL U1330 ( .A0(n1233), .A1(n386), .B0(n1247), .B1(n411), .C0(n440), 
        .C1(n385), .Y(n441) );
  CLKINVX1 U1331 ( .A(n476), .Y(n1214) );
  AOI222XL U1332 ( .A0(n1231), .A1(n386), .B0(n1249), .B1(n411), .C0(n477), 
        .C1(n385), .Y(n476) );
  CLKINVX1 U1333 ( .A(n451), .Y(n1227) );
  AOI222XL U1334 ( .A0(n1232), .A1(n382), .B0(n1251), .B1(n408), .C0(n452), 
        .C1(n380), .Y(n451) );
  CLKINVX1 U1335 ( .A(n439), .Y(n1228) );
  AOI222XL U1336 ( .A0(n1233), .A1(n382), .B0(n1247), .B1(n408), .C0(n440), 
        .C1(n380), .Y(n439) );
  OAI222XL U1337 ( .A0(n1150), .A1(n331), .B0(n329), .B1(n339), .C0(n1304), 
        .C1(n340), .Y(n774) );
  OAI222XL U1338 ( .A0(n1150), .A1(n316), .B0(n314), .B1(n341), .C0(n1298), 
        .C1(n344), .Y(n777) );
  OAI222XL U1339 ( .A0(n1150), .A1(n301), .B0(n299), .B1(n349), .C0(n1292), 
        .C1(n352), .Y(n780) );
  OAI222XL U1340 ( .A0(n1150), .A1(n286), .B0(n284), .B1(n355), .C0(n1286), 
        .C1(n358), .Y(n783) );
  OAI222XL U1341 ( .A0(n1150), .A1(n271), .B0(n269), .B1(n361), .C0(n1280), 
        .C1(n364), .Y(n786) );
  OAI222XL U1342 ( .A0(n1150), .A1(n256), .B0(n254), .B1(n367), .C0(n1274), 
        .C1(n370), .Y(n789) );
  OAI222XL U1343 ( .A0(n609), .A1(n635), .B0(n1150), .B1(n604), .C0(n1262), 
        .C1(n636), .Y(n914) );
  OA21X2 U1344 ( .A0(n1258), .A1(n1240), .B0(n1151), .Y(n627) );
  AOI2BB1X1 U1345 ( .A0N(n251), .A1N(n260), .B0(n1143), .Y(n205) );
  AOI2BB1X1 U1346 ( .A0N(n254), .A1N(n260), .B0(n1144), .Y(n206) );
  AOI2BB1X1 U1347 ( .A0N(n256), .A1N(n260), .B0(n1144), .Y(n207) );
  AOI2BB1X1 U1348 ( .A0N(n1272), .A1N(n260), .B0(n1144), .Y(n208) );
  AOI2BB1X1 U1349 ( .A0N(n266), .A1N(n275), .B0(n1144), .Y(n213) );
  AOI2BB1X1 U1350 ( .A0N(n269), .A1N(n275), .B0(n1144), .Y(n214) );
  AOI2BB1X1 U1351 ( .A0N(n271), .A1N(n275), .B0(n1144), .Y(n215) );
  AOI2BB1X1 U1352 ( .A0N(n1278), .A1N(n275), .B0(n1144), .Y(n216) );
  AOI2BB1X1 U1353 ( .A0N(n281), .A1N(n290), .B0(n1145), .Y(n221) );
  AOI2BB1X1 U1354 ( .A0N(n284), .A1N(n290), .B0(n1145), .Y(n222) );
  AOI2BB1X1 U1355 ( .A0N(n286), .A1N(n290), .B0(n1145), .Y(n223) );
  AOI2BB1X1 U1356 ( .A0N(n1284), .A1N(n290), .B0(n1145), .Y(n224) );
  AOI2BB1X1 U1357 ( .A0N(n296), .A1N(n305), .B0(n1146), .Y(n229) );
  AOI2BB1X1 U1358 ( .A0N(n299), .A1N(n305), .B0(n1145), .Y(n230) );
  AOI2BB1X1 U1359 ( .A0N(n301), .A1N(n305), .B0(n1146), .Y(n231) );
  AOI2BB1X1 U1360 ( .A0N(n1290), .A1N(n305), .B0(n1146), .Y(n232) );
  AOI2BB1X1 U1361 ( .A0N(n311), .A1N(n320), .B0(n1145), .Y(n237) );
  AOI2BB1X1 U1362 ( .A0N(n314), .A1N(n320), .B0(n1145), .Y(n238) );
  AOI2BB1X1 U1363 ( .A0N(n316), .A1N(n320), .B0(n1145), .Y(n239) );
  AOI2BB1X1 U1364 ( .A0N(n1296), .A1N(n320), .B0(n1146), .Y(n240) );
  AOI2BB1X1 U1365 ( .A0N(n326), .A1N(n335), .B0(n1146), .Y(n245) );
  AOI2BB1X1 U1366 ( .A0N(n329), .A1N(n335), .B0(n1145), .Y(n246) );
  AOI2BB1X1 U1367 ( .A0N(n331), .A1N(n335), .B0(n1146), .Y(n247) );
  AOI2BB1X1 U1368 ( .A0N(n1302), .A1N(n335), .B0(n1146), .Y(n248) );
  AOI2BB1X1 U1369 ( .A0N(n252), .A1N(n254), .B0(n1143), .Y(n202) );
  AOI2BB1X1 U1370 ( .A0N(n252), .A1N(n256), .B0(n1143), .Y(n203) );
  AOI2BB1X1 U1371 ( .A0N(n267), .A1N(n269), .B0(n1144), .Y(n210) );
  AOI2BB1X1 U1372 ( .A0N(n267), .A1N(n271), .B0(n1144), .Y(n211) );
  AOI2BB1X1 U1373 ( .A0N(n282), .A1N(n284), .B0(n1144), .Y(n218) );
  AOI2BB1X1 U1374 ( .A0N(n282), .A1N(n286), .B0(n1144), .Y(n219) );
  AOI2BB1X1 U1375 ( .A0N(n297), .A1N(n299), .B0(n1145), .Y(n226) );
  AOI2BB1X1 U1376 ( .A0N(n297), .A1N(n301), .B0(n1145), .Y(n227) );
  AOI2BB1X1 U1377 ( .A0N(n312), .A1N(n314), .B0(n1145), .Y(n234) );
  AOI2BB1X1 U1378 ( .A0N(n312), .A1N(n316), .B0(n1146), .Y(n235) );
  AOI2BB1X1 U1379 ( .A0N(n327), .A1N(n329), .B0(n1145), .Y(n242) );
  AOI2BB1X1 U1380 ( .A0N(n327), .A1N(n331), .B0(n1146), .Y(n243) );
  CLKINVX1 U1381 ( .A(N808), .Y(n1186) );
  NAND2X2 U1382 ( .A(n466), .B(n527), .Y(n502) );
  NAND2X1 U1383 ( .A(n1157), .B(n192), .Y(n631) );
  OAI22XL U1384 ( .A0(n1138), .A1(n631), .B0(n1204), .B1(n633), .Y(n913) );
  NOR2XL U1385 ( .A(n1140), .B(n1060), .Y(n633) );
  AND2X2 U1386 ( .A(n1059), .B(n404), .Y(n422) );
  AND2X2 U1387 ( .A(n1059), .B(n399), .Y(n436) );
  AND2X2 U1388 ( .A(n1059), .B(n395), .Y(n415) );
  AND2X2 U1389 ( .A(n1059), .B(n391), .Y(n413) );
  AND2X2 U1390 ( .A(n1059), .B(n387), .Y(n411) );
  AND2X2 U1391 ( .A(n1059), .B(n383), .Y(n408) );
  CLKINVX1 U1392 ( .A(n414), .Y(n1222) );
  AOI222XL U1393 ( .A0(n1235), .A1(n394), .B0(n415), .B1(n1246), .C0(n409), 
        .C1(n393), .Y(n414) );
  CLKINVX1 U1394 ( .A(n412), .Y(n1224) );
  AOI222XL U1395 ( .A0(n1235), .A1(n390), .B0(n413), .B1(n1246), .C0(n409), 
        .C1(n389), .Y(n412) );
  CLKINVX1 U1396 ( .A(n410), .Y(n1226) );
  AOI222XL U1397 ( .A0(n1235), .A1(n386), .B0(n411), .B1(n1246), .C0(n409), 
        .C1(n385), .Y(n410) );
  CLKINVX1 U1398 ( .A(n407), .Y(n1229) );
  AOI222XL U1399 ( .A0(n1235), .A1(n382), .B0(n408), .B1(n1246), .C0(n409), 
        .C1(n380), .Y(n407) );
  CLKINVX1 U1400 ( .A(n416), .Y(n1239) );
  AOI211X1 U1401 ( .A0(n1255), .A1(n417), .B0(n1149), .C0(n418), .Y(n416) );
  AND3X2 U1402 ( .A(n419), .B(n398), .C(n1257), .Y(n418) );
  AO22X1 U1403 ( .A0(n399), .A1(n1246), .B0(n420), .B1(n397), .Y(n417) );
  CLKINVX1 U1404 ( .A(n442), .Y(n1238) );
  AOI211X1 U1405 ( .A0(n1255), .A1(n443), .B0(n1149), .C0(n444), .Y(n442) );
  AND3X2 U1406 ( .A(n445), .B(n390), .C(n1257), .Y(n444) );
  AO22X1 U1407 ( .A0(n391), .A1(n1247), .B0(n446), .B1(n389), .Y(n443) );
  CLKINVX1 U1408 ( .A(n453), .Y(n1237) );
  AOI211X1 U1409 ( .A0(n1255), .A1(n454), .B0(n1149), .C0(n455), .Y(n453) );
  AND3X2 U1410 ( .A(n456), .B(n386), .C(n1257), .Y(n455) );
  AO22X1 U1411 ( .A0(n387), .A1(n1251), .B0(n457), .B1(n385), .Y(n454) );
  CLKINVX1 U1412 ( .A(n463), .Y(n1236) );
  AOI211X1 U1413 ( .A0(n1255), .A1(n464), .B0(n1149), .C0(n465), .Y(n463) );
  AND3X2 U1414 ( .A(n466), .B(n382), .C(n1257), .Y(n465) );
  AO22X1 U1415 ( .A0(n383), .A1(n1249), .B0(n467), .B1(n380), .Y(n464) );
  CLKINVX1 U1416 ( .A(n1141), .Y(n1167) );
  CLKINVX1 U1417 ( .A(n1142), .Y(n1166) );
  INVX3 U1418 ( .A(n193), .Y(n1255) );
  NAND2X1 U1419 ( .A(n1255), .B(n197), .Y(n605) );
  NOR2X1 U1420 ( .A(n559), .B(n1132), .Y(n445) );
  NAND2X1 U1421 ( .A(n1248), .B(n1263), .Y(n446) );
  NAND2X1 U1422 ( .A(n1250), .B(n1252), .Y(n467) );
  NAND2X1 U1423 ( .A(endpoint[1]), .B(n1138), .Y(n528) );
  CLKINVX1 U1424 ( .A(N1799), .Y(n1188) );
  CLKINVX1 U1425 ( .A(N1798), .Y(n1189) );
  CLKINVX1 U1426 ( .A(N1797), .Y(n1190) );
  CLKINVX1 U1427 ( .A(N1800), .Y(n1187) );
  MXI2X1 U1428 ( .A(n1095), .B(n1103), .S0(n1132), .Y(N1777) );
  MXI3X1 U1429 ( .A(n1341), .B(n1094), .C(n1095), .S0(n1117), .S1(n1121), .Y(
        N1792) );
  NAND2X1 U1430 ( .A(n258), .B(n1275), .Y(n252) );
  NAND2X1 U1431 ( .A(n273), .B(n1281), .Y(n267) );
  NAND2X1 U1432 ( .A(n288), .B(n1287), .Y(n282) );
  NAND2X1 U1433 ( .A(n303), .B(n1293), .Y(n297) );
  NAND2X1 U1434 ( .A(n318), .B(n1299), .Y(n312) );
  NAND2X1 U1435 ( .A(n333), .B(n1305), .Y(n327) );
  INVX3 U1436 ( .A(n420), .Y(n1246) );
  INVX3 U1437 ( .A(n377), .Y(n1261) );
  INVX3 U1438 ( .A(n192), .Y(n1257) );
  CLKBUFX3 U1439 ( .A(n1260), .Y(n1133) );
  CLKINVX1 U1440 ( .A(n1132), .Y(n1260) );
  OR2X1 U1441 ( .A(n1132), .B(endpoint[1]), .Y(n1067) );
  CLKBUFX3 U1442 ( .A(n1120), .Y(n1118) );
  CLKBUFX3 U1443 ( .A(endpoint[1]), .Y(n1120) );
  MXI2X1 U1444 ( .A(n1083), .B(n1097), .S0(n1121), .Y(N1783) );
  MXI3X1 U1445 ( .A(n1312), .B(n1082), .C(n1083), .S0(n1116), .S1(n1121), .Y(
        N1786) );
  CLKINVX1 U1446 ( .A(n1138), .Y(n1137) );
  INVX3 U1447 ( .A(n630), .Y(n1256) );
  CLKINVX1 U1448 ( .A(N1793), .Y(n1194) );
  CLKINVX1 U1449 ( .A(N1796), .Y(n1191) );
  CLKINVX1 U1450 ( .A(N1795), .Y(n1192) );
  NOR2X1 U1451 ( .A(n559), .B(n1133), .Y(n456) );
  NOR2X1 U1452 ( .A(n528), .B(n1132), .Y(n419) );
  CLKINVX1 U1453 ( .A(n198), .Y(n1258) );
  NAND2BX1 U1454 ( .AN(n637), .B(n638), .Y(n609) );
  NOR2X1 U1455 ( .A(n1274), .B(n1273), .Y(n369) );
  NOR2X1 U1456 ( .A(n1280), .B(n1279), .Y(n363) );
  NOR2X1 U1457 ( .A(n1286), .B(n1285), .Y(n357) );
  NOR2X1 U1458 ( .A(n1292), .B(n1291), .Y(n351) );
  NOR2X1 U1459 ( .A(n1298), .B(n1297), .Y(n343) );
  NOR2X1 U1460 ( .A(n1304), .B(n1303), .Y(n374) );
  NAND2X1 U1461 ( .A(n1274), .B(n1273), .Y(n251) );
  NAND2X1 U1462 ( .A(n1280), .B(n1279), .Y(n266) );
  NAND2X1 U1463 ( .A(n1286), .B(n1285), .Y(n281) );
  NAND2X1 U1464 ( .A(n1292), .B(n1291), .Y(n296) );
  NAND2X1 U1465 ( .A(n1298), .B(n1297), .Y(n311) );
  NAND2X1 U1466 ( .A(n1304), .B(n1303), .Y(n326) );
  AOI2BB1XL U1467 ( .A0N(num[2]), .A1N(n1062), .B0(n1245), .Y(n541) );
  AOI222XL U1468 ( .A0(\SET[3][2] ), .A1(n1267), .B0(\SET[5][2] ), .B1(n1268), 
        .C0(\SET[4][2] ), .C1(n1264), .Y(n650) );
  AOI2BB2XL U1469 ( .B0(n1124), .B1(\SET[1][2] ), .A0N(n1318), .A1N(n1062), 
        .Y(n649) );
  AOI2BB2XL U1470 ( .B0(n1124), .B1(\SET[1][4] ), .A0N(n1328), .A1N(n1062), 
        .Y(n653) );
  AOI2BB2XL U1471 ( .B0(\SET[2][2] ), .B1(n1061), .A0N(n420), .A1N(n1317), .Y(
        n665) );
  AOI222XL U1472 ( .A0(\SET[3][2] ), .A1(n1248), .B0(\SET[5][2] ), .B1(n1250), 
        .C0(\SET[4][2] ), .C1(n1064), .Y(n666) );
  AOI2BB2XL U1473 ( .B0(\SET[2][4] ), .B1(n1061), .A0N(n420), .A1N(n1327), .Y(
        n669) );
  AOI222XL U1474 ( .A0(\SET[3][4] ), .A1(n1248), .B0(\SET[5][4] ), .B1(n1250), 
        .C0(\SET[4][4] ), .C1(n1064), .Y(n670) );
  OAI221XL U1475 ( .A0(n438), .A1(n1187), .B0(n1342), .B1(n529), .C0(n530), 
        .Y(n819) );
  AOI222XL U1476 ( .A0(CNT3[7]), .A1(n1135), .B0(n531), .B1(N807), .C0(n532), 
        .C1(N821), .Y(n530) );
  OAI221XL U1477 ( .A0(n438), .A1(n1188), .B0(n1338), .B1(n529), .C0(n533), 
        .Y(n820) );
  AOI222XL U1478 ( .A0(CNT3[6]), .A1(n1135), .B0(n531), .B1(N808), .C0(n532), 
        .C1(n1125), .Y(n533) );
  OAI221XL U1479 ( .A0(n438), .A1(n1189), .B0(n1333), .B1(n529), .C0(n534), 
        .Y(n821) );
  AOI222XL U1480 ( .A0(CNT3[5]), .A1(n1135), .B0(n531), .B1(n1122), .C0(n532), 
        .C1(N823), .Y(n534) );
  OAI221XL U1481 ( .A0(n438), .A1(n1190), .B0(n1328), .B1(n529), .C0(n535), 
        .Y(n822) );
  AOI222XL U1482 ( .A0(CNT3[4]), .A1(n1135), .B0(n531), .B1(N810), .C0(n532), 
        .C1(N824), .Y(n535) );
  OAI221XL U1483 ( .A0(n438), .A1(n1191), .B0(n1323), .B1(n529), .C0(n536), 
        .Y(n823) );
  AOI222XL U1484 ( .A0(CNT3[3]), .A1(n1135), .B0(n531), .B1(n1123), .C0(n532), 
        .C1(N825), .Y(n536) );
  OAI221XL U1485 ( .A0(n438), .A1(n1192), .B0(n1318), .B1(n529), .C0(n537), 
        .Y(n824) );
  AOI222XL U1486 ( .A0(CNT3[2]), .A1(n1135), .B0(n531), .B1(N812), .C0(n532), 
        .C1(N826), .Y(n537) );
  OAI221XL U1487 ( .A0(n438), .A1(n1193), .B0(n1313), .B1(n529), .C0(n538), 
        .Y(n825) );
  AOI222XL U1488 ( .A0(CNT3[1]), .A1(n1135), .B0(n531), .B1(N813), .C0(n532), 
        .C1(N827), .Y(n538) );
  OAI221XL U1489 ( .A0(n438), .A1(n1194), .B0(n1308), .B1(n529), .C0(n539), 
        .Y(n826) );
  AOI222XL U1490 ( .A0(CNT3[0]), .A1(n1135), .B0(n531), .B1(N814), .C0(n532), 
        .C1(N828), .Y(n539) );
  CLKBUFX3 U1491 ( .A(reset), .Y(n1139) );
  NAND2X1 U1492 ( .A(n81), .B(n1138), .Y(n596) );
  OAI21XL U1493 ( .A0(n1066), .A1(n598), .B0(n1243), .Y(n597) );
  AOI2BB2XL U1494 ( .B0(\SET[2][1] ), .B1(n1061), .A0N(n420), .A1N(n1312), .Y(
        n663) );
  AOI222XL U1495 ( .A0(\SET[3][1] ), .A1(n1248), .B0(\SET[5][1] ), .B1(n1250), 
        .C0(\SET[4][1] ), .C1(n1064), .Y(n664) );
  AOI222XL U1496 ( .A0(\SET[3][1] ), .A1(n1267), .B0(\SET[5][1] ), .B1(n1268), 
        .C0(\SET[4][1] ), .C1(n1264), .Y(n648) );
  AOI2BB2XL U1497 ( .B0(n1124), .B1(\SET[1][1] ), .A0N(n1313), .A1N(n1062), 
        .Y(n647) );
  AOI222XL U1498 ( .A0(\SET[3][5] ), .A1(n1267), .B0(\SET[5][5] ), .B1(n1268), 
        .C0(\SET[4][5] ), .C1(n1264), .Y(n656) );
  AOI2BB2XL U1499 ( .B0(n1124), .B1(\SET[1][5] ), .A0N(n1333), .A1N(n1062), 
        .Y(n655) );
  AOI222XL U1500 ( .A0(\SET[3][3] ), .A1(n1267), .B0(\SET[5][3] ), .B1(n1268), 
        .C0(\SET[4][3] ), .C1(n1264), .Y(n652) );
  AOI2BB2XL U1501 ( .B0(n1124), .B1(\SET[1][3] ), .A0N(n1323), .A1N(n1062), 
        .Y(n651) );
  AOI2BB2XL U1502 ( .B0(\SET[2][0] ), .B1(n1061), .A0N(n420), .A1N(n1307), .Y(
        n661) );
  AOI222XL U1503 ( .A0(\SET[3][0] ), .A1(n1248), .B0(\SET[5][0] ), .B1(n1250), 
        .C0(\SET[4][0] ), .C1(n1064), .Y(n662) );
  AOI222XL U1504 ( .A0(\SET[3][0] ), .A1(n1267), .B0(\SET[5][0] ), .B1(n1268), 
        .C0(\SET[4][0] ), .C1(n1264), .Y(n646) );
  AOI2BB2XL U1505 ( .B0(n1124), .B1(\SET[1][0] ), .A0N(n1308), .A1N(n1062), 
        .Y(n645) );
  OAI21XL U1506 ( .A0(n445), .A1(n433), .B0(n1257), .Y(n557) );
  NAND3X1 U1507 ( .A(n1257), .B(n377), .C(n1137), .Y(n589) );
  OAI222XL U1508 ( .A0(n1230), .A1(n1193), .B0(n1196), .B1(n510), .C0(n504), 
        .C1(n89), .Y(n809) );
  AOI222XL U1509 ( .A0(CNT1[1]), .A1(n1134), .B0(n1208), .B1(N827), .C0(n1209), 
        .C1(N813), .Y(n510) );
  OAI222XL U1510 ( .A0(n1230), .A1(n1187), .B0(n1196), .B1(n595), .C0(n504), 
        .C1(n83), .Y(n852) );
  AOI222XL U1511 ( .A0(CNT1[7]), .A1(n1135), .B0(n1208), .B1(N821), .C0(n1209), 
        .C1(N807), .Y(n595) );
  OAI222XL U1512 ( .A0(n1230), .A1(n1190), .B0(n1196), .B1(n507), .C0(n504), 
        .C1(n86), .Y(n806) );
  AOI222XL U1513 ( .A0(CNT1[4]), .A1(n1134), .B0(n1208), .B1(N824), .C0(n1209), 
        .C1(N810), .Y(n507) );
  OAI222XL U1514 ( .A0(n1230), .A1(n1192), .B0(n1196), .B1(n509), .C0(n504), 
        .C1(n88), .Y(n808) );
  AOI222XL U1515 ( .A0(CNT1[2]), .A1(n1134), .B0(n1208), .B1(N826), .C0(n1209), 
        .C1(N812), .Y(n509) );
  OAI222XL U1516 ( .A0(n1230), .A1(n1188), .B0(n1196), .B1(n503), .C0(n84), 
        .C1(n504), .Y(n804) );
  AOI222XL U1517 ( .A0(CNT1[6]), .A1(n1134), .B0(n1208), .B1(n1125), .C0(n1209), .C1(N808), .Y(n503) );
  OAI222XL U1518 ( .A0(n1230), .A1(n1194), .B0(n1196), .B1(n511), .C0(n504), 
        .C1(n90), .Y(n810) );
  AOI222XL U1519 ( .A0(CNT1[0]), .A1(n1134), .B0(n1208), .B1(N828), .C0(n1209), 
        .C1(N814), .Y(n511) );
  OAI222XL U1520 ( .A0(n1230), .A1(n1189), .B0(n1196), .B1(n506), .C0(n504), 
        .C1(n85), .Y(n805) );
  AOI222XL U1521 ( .A0(CNT1[5]), .A1(n1134), .B0(n1208), .B1(N823), .C0(n1209), 
        .C1(n1122), .Y(n506) );
  OAI222XL U1522 ( .A0(n1230), .A1(n1191), .B0(n1196), .B1(n508), .C0(n504), 
        .C1(n87), .Y(n807) );
  AOI222XL U1523 ( .A0(CNT1[3]), .A1(n1134), .B0(n1208), .B1(N825), .C0(n1209), 
        .C1(n1123), .Y(n508) );
  OAI221XL U1524 ( .A0(n462), .A1(n1190), .B0(n1330), .B1(n560), .C0(n566), 
        .Y(n838) );
  CLKINVX1 U1525 ( .A(\SET[4][4] ), .Y(n1330) );
  AOI222XL U1526 ( .A0(CNT5[4]), .A1(n1136), .B0(n562), .B1(N810), .C0(n563), 
        .C1(N824), .Y(n566) );
  OAI221XL U1527 ( .A0(n450), .A1(n1190), .B0(n1329), .B1(n543), .C0(n549), 
        .Y(n830) );
  CLKINVX1 U1528 ( .A(\SET[3][4] ), .Y(n1329) );
  AOI222XL U1529 ( .A0(CNT4[4]), .A1(n1136), .B0(n545), .B1(N810), .C0(n546), 
        .C1(N824), .Y(n549) );
  OAI221XL U1530 ( .A0(n424), .A1(n1190), .B0(n1327), .B1(n512), .C0(n518), 
        .Y(n814) );
  AOI222XL U1531 ( .A0(CNT2[4]), .A1(n1134), .B0(n514), .B1(N810), .C0(n515), 
        .C1(N824), .Y(n518) );
  OAI221XL U1532 ( .A0(n502), .A1(n1190), .B0(n1326), .B1(n575), .C0(n581), 
        .Y(n846) );
  CLKINVX1 U1533 ( .A(\SET[5][4] ), .Y(n1326) );
  AOI222XL U1534 ( .A0(CNT6[4]), .A1(n505), .B0(n577), .B1(N810), .C0(n578), 
        .C1(N824), .Y(n581) );
  OAI221XL U1535 ( .A0(n462), .A1(n1192), .B0(n1320), .B1(n560), .C0(n568), 
        .Y(n840) );
  CLKINVX1 U1536 ( .A(\SET[4][2] ), .Y(n1320) );
  AOI222XL U1537 ( .A0(CNT5[2]), .A1(n1134), .B0(n562), .B1(N812), .C0(n563), 
        .C1(N826), .Y(n568) );
  OAI221XL U1538 ( .A0(n450), .A1(n1192), .B0(n1319), .B1(n543), .C0(n551), 
        .Y(n832) );
  CLKINVX1 U1539 ( .A(\SET[3][2] ), .Y(n1319) );
  AOI222XL U1540 ( .A0(CNT4[2]), .A1(n1136), .B0(n545), .B1(N812), .C0(n546), 
        .C1(N826), .Y(n551) );
  OAI221XL U1541 ( .A0(n424), .A1(n1192), .B0(n1317), .B1(n512), .C0(n520), 
        .Y(n816) );
  AOI222XL U1542 ( .A0(CNT2[2]), .A1(n1135), .B0(n514), .B1(N812), .C0(n515), 
        .C1(N826), .Y(n520) );
  OAI221XL U1543 ( .A0(n502), .A1(n1192), .B0(n1316), .B1(n575), .C0(n583), 
        .Y(n848) );
  CLKINVX1 U1544 ( .A(\SET[5][2] ), .Y(n1316) );
  AOI222XL U1545 ( .A0(CNT6[2]), .A1(n1136), .B0(n577), .B1(N812), .C0(n578), 
        .C1(N826), .Y(n583) );
  CLKBUFX3 U1546 ( .A(N811), .Y(n1123) );
  OAI211X1 U1547 ( .A0(n405), .A1(n87), .B0(n667), .C0(n668), .Y(N811) );
  AOI2BB2XL U1548 ( .B0(\SET[2][3] ), .B1(n1061), .A0N(n420), .A1N(n1322), .Y(
        n667) );
  AOI222XL U1549 ( .A0(\SET[3][3] ), .A1(n1248), .B0(\SET[5][3] ), .B1(n1250), 
        .C0(\SET[4][3] ), .C1(n1064), .Y(n668) );
  INVX3 U1550 ( .A(n615), .Y(n1199) );
  OAI31XL U1551 ( .A0(n1242), .A1(gray_data[1]), .A2(n613), .B0(n1163), .Y(
        n615) );
  INVX3 U1552 ( .A(n612), .Y(n1198) );
  OAI31XL U1553 ( .A0(n1241), .A1(gray_data[0]), .A2(n613), .B0(n1163), .Y(
        n612) );
  INVX3 U1554 ( .A(n622), .Y(n1202) );
  OAI31XL U1555 ( .A0(n618), .A1(gray_data[1]), .A2(gray_data[0]), .B0(n1163), 
        .Y(n622) );
  NOR4X1 U1556 ( .A(gray_data[3]), .B(n1258), .C(n1240), .D(n626), .Y(n623) );
  OR4X1 U1557 ( .A(gray_data[7]), .B(gray_data[6]), .C(gray_data[5]), .D(
        gray_data[4]), .Y(n626) );
  OAI221XL U1558 ( .A0(n502), .A1(n1187), .B0(n1345), .B1(n575), .C0(n576), 
        .Y(n843) );
  CLKINVX1 U1559 ( .A(\SET[5][7] ), .Y(n1345) );
  AOI222XL U1560 ( .A0(CNT6[7]), .A1(n1136), .B0(n577), .B1(N807), .C0(n578), 
        .C1(N821), .Y(n576) );
  OAI221XL U1561 ( .A0(n462), .A1(n1187), .B0(n1344), .B1(n560), .C0(n561), 
        .Y(n835) );
  CLKINVX1 U1562 ( .A(\SET[4][7] ), .Y(n1344) );
  AOI222XL U1563 ( .A0(CNT5[7]), .A1(n1136), .B0(n562), .B1(N807), .C0(n563), 
        .C1(N821), .Y(n561) );
  OAI221XL U1564 ( .A0(n450), .A1(n1187), .B0(n1343), .B1(n543), .C0(n544), 
        .Y(n827) );
  CLKINVX1 U1565 ( .A(\SET[3][7] ), .Y(n1343) );
  AOI222XL U1566 ( .A0(CNT4[7]), .A1(n1135), .B0(n545), .B1(N807), .C0(n546), 
        .C1(N821), .Y(n544) );
  OAI221XL U1567 ( .A0(n424), .A1(n1187), .B0(n1341), .B1(n512), .C0(n513), 
        .Y(n811) );
  AOI222XL U1568 ( .A0(CNT2[7]), .A1(n1134), .B0(n514), .B1(N807), .C0(n515), 
        .C1(N821), .Y(n513) );
  OAI221XL U1569 ( .A0(n462), .A1(n1188), .B0(n1340), .B1(n560), .C0(n564), 
        .Y(n836) );
  CLKINVX1 U1570 ( .A(\SET[4][6] ), .Y(n1340) );
  AOI222XL U1571 ( .A0(CNT5[6]), .A1(n1136), .B0(n562), .B1(N808), .C0(n563), 
        .C1(n1125), .Y(n564) );
  OAI221XL U1572 ( .A0(n450), .A1(n1188), .B0(n1339), .B1(n543), .C0(n547), 
        .Y(n828) );
  CLKINVX1 U1573 ( .A(\SET[3][6] ), .Y(n1339) );
  AOI222XL U1574 ( .A0(CNT4[6]), .A1(n1136), .B0(n545), .B1(N808), .C0(n546), 
        .C1(n1125), .Y(n547) );
  OAI221XL U1575 ( .A0(n424), .A1(n1188), .B0(n1337), .B1(n512), .C0(n516), 
        .Y(n812) );
  AOI222XL U1576 ( .A0(CNT2[6]), .A1(n1134), .B0(n514), .B1(N808), .C0(n515), 
        .C1(n1125), .Y(n516) );
  OAI221XL U1577 ( .A0(n502), .A1(n1188), .B0(n1336), .B1(n575), .C0(n579), 
        .Y(n844) );
  CLKINVX1 U1578 ( .A(\SET[5][6] ), .Y(n1336) );
  AOI222XL U1579 ( .A0(CNT6[6]), .A1(n1136), .B0(n577), .B1(N808), .C0(n578), 
        .C1(n1125), .Y(n579) );
  OAI221XL U1580 ( .A0(n462), .A1(n1189), .B0(n1335), .B1(n560), .C0(n565), 
        .Y(n837) );
  CLKINVX1 U1581 ( .A(\SET[4][5] ), .Y(n1335) );
  AOI222XL U1582 ( .A0(CNT5[5]), .A1(n1136), .B0(n562), .B1(n1122), .C0(n563), 
        .C1(N823), .Y(n565) );
  OAI221XL U1583 ( .A0(n450), .A1(n1189), .B0(n1334), .B1(n543), .C0(n548), 
        .Y(n829) );
  CLKINVX1 U1584 ( .A(\SET[3][5] ), .Y(n1334) );
  AOI222XL U1585 ( .A0(CNT4[5]), .A1(n1136), .B0(n545), .B1(n1122), .C0(n546), 
        .C1(N823), .Y(n548) );
  OAI221XL U1586 ( .A0(n424), .A1(n1189), .B0(n1332), .B1(n512), .C0(n517), 
        .Y(n813) );
  AOI222XL U1587 ( .A0(CNT2[5]), .A1(n1134), .B0(n514), .B1(n1122), .C0(n515), 
        .C1(N823), .Y(n517) );
  OAI221XL U1588 ( .A0(n502), .A1(n1189), .B0(n1331), .B1(n575), .C0(n580), 
        .Y(n845) );
  CLKINVX1 U1589 ( .A(\SET[5][5] ), .Y(n1331) );
  AOI222XL U1590 ( .A0(CNT6[5]), .A1(n505), .B0(n577), .B1(n1122), .C0(n578), 
        .C1(N823), .Y(n580) );
  OAI221XL U1591 ( .A0(n462), .A1(n1191), .B0(n1325), .B1(n560), .C0(n567), 
        .Y(n839) );
  CLKINVX1 U1592 ( .A(\SET[4][3] ), .Y(n1325) );
  AOI222XL U1593 ( .A0(CNT5[3]), .A1(n1136), .B0(n562), .B1(n1123), .C0(n563), 
        .C1(N825), .Y(n567) );
  OAI221XL U1594 ( .A0(n450), .A1(n1191), .B0(n1324), .B1(n543), .C0(n550), 
        .Y(n831) );
  CLKINVX1 U1595 ( .A(\SET[3][3] ), .Y(n1324) );
  AOI222XL U1596 ( .A0(CNT4[3]), .A1(n1136), .B0(n545), .B1(n1123), .C0(n546), 
        .C1(N825), .Y(n550) );
  OAI221XL U1597 ( .A0(n424), .A1(n1191), .B0(n1322), .B1(n512), .C0(n519), 
        .Y(n815) );
  AOI222XL U1598 ( .A0(CNT2[3]), .A1(n1134), .B0(n514), .B1(n1123), .C0(n515), 
        .C1(N825), .Y(n519) );
  OAI221XL U1599 ( .A0(n502), .A1(n1191), .B0(n1321), .B1(n575), .C0(n582), 
        .Y(n847) );
  CLKINVX1 U1600 ( .A(\SET[5][3] ), .Y(n1321) );
  AOI222XL U1601 ( .A0(CNT6[3]), .A1(n1135), .B0(n577), .B1(n1123), .C0(n578), 
        .C1(N825), .Y(n582) );
  OAI221XL U1602 ( .A0(n462), .A1(n1193), .B0(n1315), .B1(n560), .C0(n569), 
        .Y(n841) );
  CLKINVX1 U1603 ( .A(\SET[4][1] ), .Y(n1315) );
  AOI222XL U1604 ( .A0(CNT5[1]), .A1(n1134), .B0(n562), .B1(N813), .C0(n563), 
        .C1(N827), .Y(n569) );
  OAI221XL U1605 ( .A0(n450), .A1(n1193), .B0(n1314), .B1(n543), .C0(n552), 
        .Y(n833) );
  CLKINVX1 U1606 ( .A(\SET[3][1] ), .Y(n1314) );
  AOI222XL U1607 ( .A0(CNT4[1]), .A1(n1136), .B0(n545), .B1(N813), .C0(n546), 
        .C1(N827), .Y(n552) );
  OAI221XL U1608 ( .A0(n424), .A1(n1193), .B0(n1312), .B1(n512), .C0(n521), 
        .Y(n817) );
  AOI222XL U1609 ( .A0(CNT2[1]), .A1(n1135), .B0(n514), .B1(N813), .C0(n515), 
        .C1(N827), .Y(n521) );
  OAI221XL U1610 ( .A0(n502), .A1(n1193), .B0(n1311), .B1(n575), .C0(n584), 
        .Y(n849) );
  CLKINVX1 U1611 ( .A(\SET[5][1] ), .Y(n1311) );
  AOI222XL U1612 ( .A0(CNT6[1]), .A1(n1136), .B0(n577), .B1(N813), .C0(n578), 
        .C1(N827), .Y(n584) );
  OAI221XL U1613 ( .A0(n462), .A1(n1194), .B0(n1310), .B1(n560), .C0(n570), 
        .Y(n842) );
  CLKINVX1 U1614 ( .A(\SET[4][0] ), .Y(n1310) );
  AOI222XL U1615 ( .A0(CNT5[0]), .A1(n1135), .B0(n562), .B1(N814), .C0(n563), 
        .C1(N828), .Y(n570) );
  OAI221XL U1616 ( .A0(n450), .A1(n1194), .B0(n1309), .B1(n543), .C0(n553), 
        .Y(n834) );
  CLKINVX1 U1617 ( .A(\SET[3][0] ), .Y(n1309) );
  AOI222XL U1618 ( .A0(CNT4[0]), .A1(n1136), .B0(n545), .B1(N814), .C0(n546), 
        .C1(N828), .Y(n553) );
  OAI221XL U1619 ( .A0(n424), .A1(n1194), .B0(n1307), .B1(n512), .C0(n522), 
        .Y(n818) );
  AOI222XL U1620 ( .A0(CNT2[0]), .A1(n1135), .B0(n514), .B1(N814), .C0(n515), 
        .C1(N828), .Y(n522) );
  OAI221XL U1621 ( .A0(n502), .A1(n1194), .B0(n1306), .B1(n575), .C0(n585), 
        .Y(n850) );
  CLKINVX1 U1622 ( .A(\SET[5][0] ), .Y(n1306) );
  AOI222XL U1623 ( .A0(CNT6[0]), .A1(n1134), .B0(n577), .B1(N814), .C0(n578), 
        .C1(N828), .Y(n585) );
  INVX3 U1624 ( .A(n620), .Y(n1201) );
  OAI31XL U1625 ( .A0(n618), .A1(gray_data[1]), .A2(n1242), .B0(n1160), .Y(
        n620) );
  INVX3 U1626 ( .A(n617), .Y(n1200) );
  OAI31XL U1627 ( .A0(n618), .A1(gray_data[0]), .A2(n1241), .B0(n1159), .Y(
        n617) );
  NAND2X1 U1628 ( .A(num[1]), .B(num[0]), .Y(n558) );
  NAND2X1 U1629 ( .A(num[2]), .B(num[0]), .Y(n590) );
  NAND2X1 U1630 ( .A(num[2]), .B(n1265), .Y(n574) );
  NAND2BX1 U1631 ( .AN(gray_data[2]), .B(n623), .Y(n613) );
  NAND2X1 U1632 ( .A(gray_data[2]), .B(n623), .Y(n618) );
  CLKBUFX3 U1633 ( .A(n474), .Y(n1124) );
  CLKINVX1 U1634 ( .A(\SET[1][2] ), .Y(n1317) );
  CLKINVX1 U1635 ( .A(\SET[1][1] ), .Y(n1312) );
  CLKINVX1 U1636 ( .A(\SET[1][4] ), .Y(n1327) );
  CLKINVX1 U1637 ( .A(\SET[2][1] ), .Y(n1313) );
  CLKINVX1 U1638 ( .A(\SET[2][2] ), .Y(n1318) );
  CLKINVX1 U1639 ( .A(\SET[2][5] ), .Y(n1333) );
  CLKINVX1 U1640 ( .A(\SET[2][4] ), .Y(n1328) );
  CLKINVX1 U1641 ( .A(\SET[2][3] ), .Y(n1323) );
  AO22X1 U1642 ( .A0(n1203), .A1(CNT3[0]), .B0(N908), .B1(n624), .Y(n902) );
  AO22X1 U1643 ( .A0(n1199), .A1(CNT1[0]), .B0(N892), .B1(n614), .Y(n870) );
  AO22X1 U1644 ( .A0(n1198), .A1(CNT2[0]), .B0(N900), .B1(n611), .Y(n862) );
  AO22X1 U1645 ( .A0(n1202), .A1(CNT4[0]), .B0(N916), .B1(n621), .Y(n894) );
  AO22X1 U1646 ( .A0(n1201), .A1(CNT5[0]), .B0(N924), .B1(n619), .Y(n886) );
  AO22X1 U1647 ( .A0(n1200), .A1(CNT6[0]), .B0(N932), .B1(n616), .Y(n878) );
  AO22X1 U1648 ( .A0(n1203), .A1(CNT3[6]), .B0(N914), .B1(n624), .Y(n896) );
  AO22X1 U1649 ( .A0(n1203), .A1(CNT3[5]), .B0(N913), .B1(n624), .Y(n897) );
  AO22X1 U1650 ( .A0(n1203), .A1(CNT3[4]), .B0(N912), .B1(n624), .Y(n898) );
  AO22X1 U1651 ( .A0(n1203), .A1(CNT3[3]), .B0(N911), .B1(n624), .Y(n899) );
  AO22X1 U1652 ( .A0(n1203), .A1(CNT3[2]), .B0(N910), .B1(n624), .Y(n900) );
  AO22X1 U1653 ( .A0(n1203), .A1(CNT3[1]), .B0(N909), .B1(n624), .Y(n901) );
  AO22X1 U1654 ( .A0(n1199), .A1(CNT1[6]), .B0(N898), .B1(n614), .Y(n864) );
  AO22X1 U1655 ( .A0(n1199), .A1(CNT1[5]), .B0(N897), .B1(n614), .Y(n865) );
  AO22X1 U1656 ( .A0(n1199), .A1(CNT1[4]), .B0(N896), .B1(n614), .Y(n866) );
  AO22X1 U1657 ( .A0(n1199), .A1(CNT1[3]), .B0(N895), .B1(n614), .Y(n867) );
  AO22X1 U1658 ( .A0(n1199), .A1(CNT1[2]), .B0(N894), .B1(n614), .Y(n868) );
  AO22X1 U1659 ( .A0(n1199), .A1(CNT1[1]), .B0(N893), .B1(n614), .Y(n869) );
  AO22X1 U1660 ( .A0(n1198), .A1(CNT2[6]), .B0(N906), .B1(n611), .Y(n856) );
  AO22X1 U1661 ( .A0(n1198), .A1(CNT2[5]), .B0(N905), .B1(n611), .Y(n857) );
  AO22X1 U1662 ( .A0(n1198), .A1(CNT2[4]), .B0(N904), .B1(n611), .Y(n858) );
  AO22X1 U1663 ( .A0(n1198), .A1(CNT2[3]), .B0(N903), .B1(n611), .Y(n859) );
  AO22X1 U1664 ( .A0(n1198), .A1(CNT2[2]), .B0(N902), .B1(n611), .Y(n860) );
  AO22X1 U1665 ( .A0(n1198), .A1(CNT2[1]), .B0(N901), .B1(n611), .Y(n861) );
  AO22X1 U1666 ( .A0(n1202), .A1(CNT4[6]), .B0(N922), .B1(n621), .Y(n888) );
  AO22X1 U1667 ( .A0(n1202), .A1(CNT4[5]), .B0(N921), .B1(n621), .Y(n889) );
  AO22X1 U1668 ( .A0(n1202), .A1(CNT4[4]), .B0(N920), .B1(n621), .Y(n890) );
  AO22X1 U1669 ( .A0(n1202), .A1(CNT4[3]), .B0(N919), .B1(n621), .Y(n891) );
  AO22X1 U1670 ( .A0(n1202), .A1(CNT4[2]), .B0(N918), .B1(n621), .Y(n892) );
  AO22X1 U1671 ( .A0(n1202), .A1(CNT4[1]), .B0(N917), .B1(n621), .Y(n893) );
  AO22X1 U1672 ( .A0(n1201), .A1(CNT5[6]), .B0(N930), .B1(n619), .Y(n880) );
  AO22X1 U1673 ( .A0(n1201), .A1(CNT5[5]), .B0(N929), .B1(n619), .Y(n881) );
  AO22X1 U1674 ( .A0(n1201), .A1(CNT5[4]), .B0(N928), .B1(n619), .Y(n882) );
  AO22X1 U1675 ( .A0(n1201), .A1(CNT5[3]), .B0(N927), .B1(n619), .Y(n883) );
  AO22X1 U1676 ( .A0(n1201), .A1(CNT5[2]), .B0(N926), .B1(n619), .Y(n884) );
  AO22X1 U1677 ( .A0(n1201), .A1(CNT5[1]), .B0(N925), .B1(n619), .Y(n885) );
  AO22X1 U1678 ( .A0(n1200), .A1(CNT6[6]), .B0(N938), .B1(n616), .Y(n872) );
  AO22X1 U1679 ( .A0(n1200), .A1(CNT6[5]), .B0(N937), .B1(n616), .Y(n873) );
  AO22X1 U1680 ( .A0(n1200), .A1(CNT6[4]), .B0(N936), .B1(n616), .Y(n874) );
  AO22X1 U1681 ( .A0(n1200), .A1(CNT6[3]), .B0(N935), .B1(n616), .Y(n875) );
  AO22X1 U1682 ( .A0(n1200), .A1(CNT6[2]), .B0(N934), .B1(n616), .Y(n876) );
  AO22X1 U1683 ( .A0(n1200), .A1(CNT6[1]), .B0(N933), .B1(n616), .Y(n877) );
  AO22X1 U1684 ( .A0(n1203), .A1(CNT3[7]), .B0(N915), .B1(n624), .Y(n903) );
  AO22X1 U1685 ( .A0(n1199), .A1(CNT1[7]), .B0(N899), .B1(n614), .Y(n871) );
  AO22X1 U1686 ( .A0(n1198), .A1(CNT2[7]), .B0(N907), .B1(n611), .Y(n863) );
  AO22X1 U1687 ( .A0(n1202), .A1(CNT4[7]), .B0(N923), .B1(n621), .Y(n895) );
  AO22X1 U1688 ( .A0(n1201), .A1(CNT5[7]), .B0(N931), .B1(n619), .Y(n887) );
  AO22X1 U1689 ( .A0(n1200), .A1(CNT6[7]), .B0(N939), .B1(n616), .Y(n879) );
  CLKBUFX3 U1690 ( .A(N809), .Y(n1122) );
  OAI211X1 U1691 ( .A0(n405), .A1(n85), .B0(n671), .C0(n672), .Y(N809) );
  AOI2BB2X1 U1692 ( .B0(\SET[2][5] ), .B1(n1061), .A0N(n420), .A1N(n1332), .Y(
        n671) );
  AOI222XL U1693 ( .A0(\SET[3][5] ), .A1(n1248), .B0(\SET[5][5] ), .B1(n1250), 
        .C0(\SET[4][5] ), .C1(n1064), .Y(n672) );
  AOI222XL U1694 ( .A0(\SET[3][7] ), .A1(n1248), .B0(\SET[5][7] ), .B1(n1250), 
        .C0(\SET[4][7] ), .C1(n1064), .Y(n676) );
  AOI222XL U1695 ( .A0(\SET[3][6] ), .A1(n1248), .B0(\SET[5][6] ), .B1(n1250), 
        .C0(\SET[4][6] ), .C1(n1064), .Y(n674) );
  AOI222XL U1696 ( .A0(\SET[3][7] ), .A1(n1267), .B0(\SET[5][7] ), .B1(n1268), 
        .C0(\SET[4][7] ), .C1(n1264), .Y(n660) );
  OAI32X1 U1697 ( .A0(n339), .A1(\bitpos[0][2] ), .A2(n1302), .B0(n373), .B1(
        n1305), .Y(n791) );
  OA21XL U1698 ( .A0(n1150), .A1(n374), .B0(n340), .Y(n373) );
  OAI32X1 U1699 ( .A0(n341), .A1(\bitpos[1][2] ), .A2(n1296), .B0(n342), .B1(
        n1299), .Y(n776) );
  OA21XL U1700 ( .A0(n1150), .A1(n343), .B0(n344), .Y(n342) );
  OAI32X1 U1701 ( .A0(n349), .A1(\bitpos[2][2] ), .A2(n1290), .B0(n350), .B1(
        n1293), .Y(n779) );
  OA21XL U1702 ( .A0(n1150), .A1(n351), .B0(n352), .Y(n350) );
  OAI32X1 U1703 ( .A0(n355), .A1(\bitpos[3][2] ), .A2(n1284), .B0(n356), .B1(
        n1287), .Y(n782) );
  OA21XL U1704 ( .A0(n1150), .A1(n357), .B0(n358), .Y(n356) );
  OAI32X1 U1705 ( .A0(n361), .A1(\bitpos[4][2] ), .A2(n1278), .B0(n362), .B1(
        n1281), .Y(n785) );
  OA21XL U1706 ( .A0(n1150), .A1(n363), .B0(n364), .Y(n362) );
  OAI32X1 U1707 ( .A0(n367), .A1(\bitpos[5][2] ), .A2(n1272), .B0(n368), .B1(
        n1275), .Y(n788) );
  OA21XL U1708 ( .A0(n1150), .A1(n369), .B0(n370), .Y(n368) );
  OAI31XL U1709 ( .A0(n199), .A1(state[0]), .A2(n1146), .B0(n200), .Y(n677) );
  NAND2X1 U1710 ( .A(code_valid), .B(n199), .Y(n200) );
  AOI2BB1X1 U1711 ( .A0N(state[1]), .A1N(n68), .B0(n1143), .Y(n199) );
  OAI31XL U1712 ( .A0(n1127), .A1(n1148), .A2(n201), .B0(n250), .Y(n726) );
  NAND2X1 U1713 ( .A(HC6[0]), .B(n201), .Y(n250) );
  OAI31XL U1714 ( .A0(n1127), .A1(n1148), .A2(n202), .B0(n253), .Y(n727) );
  NAND2X1 U1715 ( .A(HC6[1]), .B(n202), .Y(n253) );
  OAI31XL U1716 ( .A0(n1127), .A1(n1148), .A2(n203), .B0(n255), .Y(n728) );
  NAND2X1 U1717 ( .A(HC6[2]), .B(n203), .Y(n255) );
  OAI31XL U1718 ( .A0(n1127), .A1(n1149), .A2(n204), .B0(n257), .Y(n729) );
  NAND2X1 U1719 ( .A(HC6[3]), .B(n204), .Y(n257) );
  OAI31XL U1720 ( .A0(n1127), .A1(n1147), .A2(n205), .B0(n259), .Y(n730) );
  NAND2X1 U1721 ( .A(HC6[4]), .B(n205), .Y(n259) );
  OAI31XL U1722 ( .A0(n1127), .A1(n1148), .A2(n206), .B0(n261), .Y(n731) );
  NAND2X1 U1723 ( .A(HC6[5]), .B(n206), .Y(n261) );
  OAI31XL U1724 ( .A0(n1127), .A1(n1147), .A2(n207), .B0(n262), .Y(n732) );
  NAND2X1 U1725 ( .A(HC6[6]), .B(n207), .Y(n262) );
  OAI31XL U1726 ( .A0(n1127), .A1(n1149), .A2(n208), .B0(n263), .Y(n733) );
  NAND2X1 U1727 ( .A(HC6[7]), .B(n208), .Y(n263) );
  OAI31XL U1728 ( .A0(n1128), .A1(n1148), .A2(n209), .B0(n265), .Y(n734) );
  NAND2X1 U1729 ( .A(HC5[0]), .B(n209), .Y(n265) );
  OAI31XL U1730 ( .A0(n1128), .A1(n1147), .A2(n210), .B0(n268), .Y(n735) );
  NAND2X1 U1731 ( .A(HC5[1]), .B(n210), .Y(n268) );
  OAI31XL U1732 ( .A0(n1128), .A1(n1147), .A2(n211), .B0(n270), .Y(n736) );
  NAND2X1 U1733 ( .A(HC5[2]), .B(n211), .Y(n270) );
  OAI31XL U1734 ( .A0(n1128), .A1(n1148), .A2(n212), .B0(n272), .Y(n737) );
  NAND2X1 U1735 ( .A(HC5[3]), .B(n212), .Y(n272) );
  OAI31XL U1736 ( .A0(n1128), .A1(n1147), .A2(n213), .B0(n274), .Y(n738) );
  NAND2X1 U1737 ( .A(HC5[4]), .B(n213), .Y(n274) );
  OAI31XL U1738 ( .A0(n1128), .A1(n1148), .A2(n214), .B0(n276), .Y(n739) );
  NAND2X1 U1739 ( .A(HC5[5]), .B(n214), .Y(n276) );
  OAI31XL U1740 ( .A0(n1128), .A1(n1147), .A2(n215), .B0(n277), .Y(n740) );
  NAND2X1 U1741 ( .A(HC5[6]), .B(n215), .Y(n277) );
  OAI31XL U1742 ( .A0(n1128), .A1(n1148), .A2(n216), .B0(n278), .Y(n741) );
  NAND2X1 U1743 ( .A(HC5[7]), .B(n216), .Y(n278) );
  OAI31XL U1744 ( .A0(n1129), .A1(n1147), .A2(n217), .B0(n280), .Y(n742) );
  NAND2X1 U1745 ( .A(HC4[0]), .B(n217), .Y(n280) );
  OAI31XL U1746 ( .A0(n1129), .A1(n1148), .A2(n218), .B0(n283), .Y(n743) );
  NAND2X1 U1747 ( .A(HC4[1]), .B(n218), .Y(n283) );
  OAI31XL U1748 ( .A0(n1129), .A1(n1147), .A2(n219), .B0(n285), .Y(n744) );
  NAND2X1 U1749 ( .A(HC4[2]), .B(n219), .Y(n285) );
  OAI31XL U1750 ( .A0(n1129), .A1(n1148), .A2(n220), .B0(n287), .Y(n745) );
  NAND2X1 U1751 ( .A(HC4[3]), .B(n220), .Y(n287) );
  OAI31XL U1752 ( .A0(n1129), .A1(n1147), .A2(n221), .B0(n289), .Y(n746) );
  NAND2X1 U1753 ( .A(HC4[4]), .B(n221), .Y(n289) );
  OAI31XL U1754 ( .A0(n1129), .A1(n1146), .A2(n222), .B0(n291), .Y(n747) );
  NAND2X1 U1755 ( .A(HC4[5]), .B(n222), .Y(n291) );
  OAI31XL U1756 ( .A0(n1129), .A1(n1147), .A2(n223), .B0(n292), .Y(n748) );
  NAND2X1 U1757 ( .A(HC4[6]), .B(n223), .Y(n292) );
  OAI31XL U1758 ( .A0(n1129), .A1(n1147), .A2(n224), .B0(n293), .Y(n749) );
  NAND2X1 U1759 ( .A(HC4[7]), .B(n224), .Y(n293) );
  OAI31XL U1760 ( .A0(n1130), .A1(n1147), .A2(n225), .B0(n295), .Y(n750) );
  NAND2X1 U1761 ( .A(HC3[0]), .B(n225), .Y(n295) );
  OAI31XL U1762 ( .A0(n1130), .A1(n1147), .A2(n226), .B0(n298), .Y(n751) );
  NAND2X1 U1763 ( .A(HC3[1]), .B(n226), .Y(n298) );
  OAI31XL U1764 ( .A0(n1130), .A1(n1147), .A2(n227), .B0(n300), .Y(n752) );
  NAND2X1 U1765 ( .A(HC3[2]), .B(n227), .Y(n300) );
  OAI31XL U1766 ( .A0(n1130), .A1(n1147), .A2(n228), .B0(n302), .Y(n753) );
  NAND2X1 U1767 ( .A(HC3[3]), .B(n228), .Y(n302) );
  OAI31XL U1768 ( .A0(n1130), .A1(n1147), .A2(n229), .B0(n304), .Y(n754) );
  NAND2X1 U1769 ( .A(HC3[4]), .B(n229), .Y(n304) );
  OAI31XL U1770 ( .A0(n1130), .A1(n1147), .A2(n230), .B0(n306), .Y(n755) );
  NAND2X1 U1771 ( .A(HC3[5]), .B(n230), .Y(n306) );
  OAI31XL U1772 ( .A0(n1130), .A1(n1147), .A2(n231), .B0(n307), .Y(n756) );
  NAND2X1 U1773 ( .A(HC3[6]), .B(n231), .Y(n307) );
  OAI31XL U1774 ( .A0(n1130), .A1(n1148), .A2(n232), .B0(n308), .Y(n757) );
  NAND2X1 U1775 ( .A(HC3[7]), .B(n232), .Y(n308) );
  OAI31XL U1776 ( .A0(n1131), .A1(n1148), .A2(n233), .B0(n310), .Y(n758) );
  NAND2X1 U1777 ( .A(HC2[0]), .B(n233), .Y(n310) );
  OAI31XL U1778 ( .A0(n1131), .A1(n1148), .A2(n234), .B0(n313), .Y(n759) );
  NAND2X1 U1779 ( .A(HC2[1]), .B(n234), .Y(n313) );
  OAI31XL U1780 ( .A0(n1131), .A1(n1148), .A2(n235), .B0(n315), .Y(n760) );
  NAND2X1 U1781 ( .A(HC2[2]), .B(n235), .Y(n315) );
  OAI31XL U1782 ( .A0(n1131), .A1(n1148), .A2(n236), .B0(n317), .Y(n761) );
  NAND2X1 U1783 ( .A(HC2[3]), .B(n236), .Y(n317) );
  OAI31XL U1784 ( .A0(n1131), .A1(n1148), .A2(n237), .B0(n319), .Y(n762) );
  NAND2X1 U1785 ( .A(HC2[4]), .B(n237), .Y(n319) );
  OAI31XL U1786 ( .A0(n1131), .A1(n1148), .A2(n238), .B0(n321), .Y(n763) );
  NAND2X1 U1787 ( .A(HC2[5]), .B(n238), .Y(n321) );
  OAI31XL U1788 ( .A0(n1131), .A1(n1149), .A2(n239), .B0(n322), .Y(n764) );
  NAND2X1 U1789 ( .A(HC2[6]), .B(n239), .Y(n322) );
  OAI31XL U1790 ( .A0(n1131), .A1(n1148), .A2(n240), .B0(n323), .Y(n765) );
  NAND2X1 U1791 ( .A(HC2[7]), .B(n240), .Y(n323) );
  OAI31XL U1792 ( .A0(n1126), .A1(n1149), .A2(n241), .B0(n325), .Y(n766) );
  NAND2X1 U1793 ( .A(HC1[0]), .B(n241), .Y(n325) );
  OAI31XL U1794 ( .A0(n1126), .A1(n1149), .A2(n242), .B0(n328), .Y(n767) );
  NAND2X1 U1795 ( .A(HC1[1]), .B(n242), .Y(n328) );
  OAI31XL U1796 ( .A0(n1126), .A1(n1149), .A2(n243), .B0(n330), .Y(n768) );
  NAND2X1 U1797 ( .A(HC1[2]), .B(n243), .Y(n330) );
  OAI31XL U1798 ( .A0(n1126), .A1(n1149), .A2(n244), .B0(n332), .Y(n769) );
  NAND2X1 U1799 ( .A(HC1[3]), .B(n244), .Y(n332) );
  OAI31XL U1800 ( .A0(n1126), .A1(n1149), .A2(n245), .B0(n334), .Y(n770) );
  NAND2X1 U1801 ( .A(HC1[4]), .B(n245), .Y(n334) );
  OAI31XL U1802 ( .A0(n1126), .A1(n1149), .A2(n246), .B0(n336), .Y(n771) );
  NAND2X1 U1803 ( .A(HC1[5]), .B(n246), .Y(n336) );
  OAI31XL U1804 ( .A0(n1126), .A1(n1149), .A2(n247), .B0(n337), .Y(n772) );
  NAND2X1 U1805 ( .A(HC1[6]), .B(n247), .Y(n337) );
  OAI31XL U1806 ( .A0(n1126), .A1(n1149), .A2(n248), .B0(n338), .Y(n773) );
  NAND2X1 U1807 ( .A(HC1[7]), .B(n248), .Y(n338) );
  OAI22XL U1808 ( .A0(n1253), .A1(n636), .B0(times[0]), .B1(n635), .Y(n915) );
  OAI22XL U1809 ( .A0(n1252), .A1(n606), .B0(n1207), .B1(n607), .Y(n855) );
  AOI22X1 U1810 ( .A0(n1209), .A1(n608), .B0(n609), .B1(n1208), .Y(n607) );
  OAI21XL U1811 ( .A0(count[1]), .A1(count[0]), .B0(n610), .Y(n608) );
  OAI22XL U1812 ( .A0(n1303), .A1(n340), .B0(\bitpos[0][0] ), .B1(n339), .Y(
        n775) );
  OAI22XL U1813 ( .A0(n1297), .A1(n344), .B0(\bitpos[1][0] ), .B1(n341), .Y(
        n778) );
  OAI22XL U1814 ( .A0(n1291), .A1(n352), .B0(\bitpos[2][0] ), .B1(n349), .Y(
        n781) );
  OAI22XL U1815 ( .A0(n1285), .A1(n358), .B0(\bitpos[3][0] ), .B1(n355), .Y(
        n784) );
  OAI22XL U1816 ( .A0(n1279), .A1(n364), .B0(\bitpos[4][0] ), .B1(n361), .Y(
        n787) );
  OAI22XL U1817 ( .A0(n1273), .A1(n370), .B0(\bitpos[5][0] ), .B1(n367), .Y(
        n790) );
  OAI22XL U1818 ( .A0(n1244), .A1(n606), .B0(n1207), .B1(n644), .Y(n918) );
  OAI22XL U1819 ( .A0(n1269), .A1(n591), .B0(n1205), .B1(n592), .Y(n851) );
  AOI2BB2X1 U1820 ( .B0(n1209), .B1(n593), .A0N(n1262), .A1N(n594), .Y(n592)
         );
  OAI21XL U1821 ( .A0(num[1]), .A1(num[0]), .B0(n558), .Y(n593) );
  OAI22XL U1822 ( .A0(n1263), .A1(n606), .B0(n1207), .B1(n640), .Y(n917) );
  AOI2BB2X1 U1823 ( .B0(n1209), .B1(n641), .A0N(n642), .A1N(n594), .Y(n640) );
  XNOR2X1 U1824 ( .A(times[2]), .B(n637), .Y(n642) );
  OAI21XL U1825 ( .A0(n1263), .A1(n1252), .B0(n643), .Y(n641) );
  AO22X1 U1826 ( .A0(n599), .A1(n591), .B0(num[2]), .B1(n600), .Y(n853) );
  OAI2BB2XL U1827 ( .B0(n602), .B1(n601), .A0N(times[2]), .A1N(n1208), .Y(n599) );
  OAI21XL U1828 ( .A0(n1269), .A1(n601), .B0(n591), .Y(n600) );
  NOR2X1 U1829 ( .A(n1268), .B(n598), .Y(n602) );
  OAI21XL U1830 ( .A0(n638), .A1(n635), .B0(n639), .Y(n916) );
  OAI21XL U1831 ( .A0(n1059), .A1(n1206), .B0(times[2]), .Y(n639) );
  OAI2BB2XL U1832 ( .B0(n1140), .B1(n201), .A0N(M6[0]), .A1N(n201), .Y(n678)
         );
  OAI2BB2XL U1833 ( .B0(n1141), .B1(n202), .A0N(M6[1]), .A1N(n202), .Y(n679)
         );
  OAI2BB2XL U1834 ( .B0(n1141), .B1(n203), .A0N(M6[2]), .A1N(n203), .Y(n680)
         );
  OAI2BB2XL U1835 ( .B0(n1141), .B1(n204), .A0N(M6[3]), .A1N(n204), .Y(n681)
         );
  OAI2BB2XL U1836 ( .B0(n1141), .B1(n205), .A0N(M6[4]), .A1N(n205), .Y(n682)
         );
  OAI2BB2XL U1837 ( .B0(n1141), .B1(n206), .A0N(M6[5]), .A1N(n206), .Y(n683)
         );
  OAI2BB2XL U1838 ( .B0(n1141), .B1(n207), .A0N(M6[6]), .A1N(n207), .Y(n684)
         );
  OAI2BB2XL U1839 ( .B0(n1141), .B1(n208), .A0N(M6[7]), .A1N(n208), .Y(n685)
         );
  OAI2BB2XL U1840 ( .B0(n1141), .B1(n209), .A0N(M5[0]), .A1N(n209), .Y(n686)
         );
  OAI2BB2XL U1841 ( .B0(n1141), .B1(n210), .A0N(M5[1]), .A1N(n210), .Y(n687)
         );
  OAI2BB2XL U1842 ( .B0(n1141), .B1(n211), .A0N(M5[2]), .A1N(n211), .Y(n688)
         );
  OAI2BB2XL U1843 ( .B0(n1141), .B1(n212), .A0N(M5[3]), .A1N(n212), .Y(n689)
         );
  OAI2BB2XL U1844 ( .B0(n1141), .B1(n213), .A0N(M5[4]), .A1N(n213), .Y(n690)
         );
  OAI2BB2XL U1845 ( .B0(n1142), .B1(n214), .A0N(M5[5]), .A1N(n214), .Y(n691)
         );
  OAI2BB2XL U1846 ( .B0(n1142), .B1(n215), .A0N(M5[6]), .A1N(n215), .Y(n692)
         );
  OAI2BB2XL U1847 ( .B0(n1141), .B1(n216), .A0N(M5[7]), .A1N(n216), .Y(n693)
         );
  OAI2BB2XL U1848 ( .B0(n1142), .B1(n217), .A0N(M4[0]), .A1N(n217), .Y(n694)
         );
  OAI2BB2XL U1849 ( .B0(n1142), .B1(n218), .A0N(M4[1]), .A1N(n218), .Y(n695)
         );
  OAI2BB2XL U1850 ( .B0(n1142), .B1(n219), .A0N(M4[2]), .A1N(n219), .Y(n696)
         );
  OAI2BB2XL U1851 ( .B0(n1142), .B1(n220), .A0N(M4[3]), .A1N(n220), .Y(n697)
         );
  OAI2BB2XL U1852 ( .B0(n1142), .B1(n221), .A0N(M4[4]), .A1N(n221), .Y(n698)
         );
  OAI2BB2XL U1853 ( .B0(n1142), .B1(n222), .A0N(M4[5]), .A1N(n222), .Y(n699)
         );
  OAI2BB2XL U1854 ( .B0(n1142), .B1(n223), .A0N(M4[6]), .A1N(n223), .Y(n700)
         );
  OAI2BB2XL U1855 ( .B0(n1142), .B1(n224), .A0N(M4[7]), .A1N(n224), .Y(n701)
         );
  OAI2BB2XL U1856 ( .B0(n1142), .B1(n225), .A0N(M3[0]), .A1N(n225), .Y(n702)
         );
  OAI2BB2XL U1857 ( .B0(n1142), .B1(n226), .A0N(M3[1]), .A1N(n226), .Y(n703)
         );
  OAI2BB2XL U1858 ( .B0(n1141), .B1(n227), .A0N(M3[2]), .A1N(n227), .Y(n704)
         );
  OAI2BB2XL U1859 ( .B0(n1142), .B1(n228), .A0N(M3[3]), .A1N(n228), .Y(n705)
         );
  OAI2BB2XL U1860 ( .B0(n1142), .B1(n229), .A0N(M3[4]), .A1N(n229), .Y(n706)
         );
  OAI2BB2XL U1861 ( .B0(n1142), .B1(n230), .A0N(M3[5]), .A1N(n230), .Y(n707)
         );
  OAI2BB2XL U1862 ( .B0(n1141), .B1(n231), .A0N(M3[6]), .A1N(n231), .Y(n708)
         );
  OAI2BB2XL U1863 ( .B0(n1142), .B1(n232), .A0N(M3[7]), .A1N(n232), .Y(n709)
         );
  OAI2BB2XL U1864 ( .B0(n1141), .B1(n233), .A0N(M2[0]), .A1N(n233), .Y(n710)
         );
  OAI2BB2XL U1865 ( .B0(n1142), .B1(n234), .A0N(M2[1]), .A1N(n234), .Y(n711)
         );
  OAI2BB2XL U1866 ( .B0(n1141), .B1(n235), .A0N(M2[2]), .A1N(n235), .Y(n712)
         );
  OAI2BB2XL U1867 ( .B0(n1142), .B1(n236), .A0N(M2[3]), .A1N(n236), .Y(n713)
         );
  OAI2BB2XL U1868 ( .B0(n1141), .B1(n237), .A0N(M2[4]), .A1N(n237), .Y(n714)
         );
  OAI2BB2XL U1869 ( .B0(n1142), .B1(n238), .A0N(M2[5]), .A1N(n238), .Y(n715)
         );
  OAI2BB2XL U1870 ( .B0(n1141), .B1(n239), .A0N(M2[6]), .A1N(n239), .Y(n716)
         );
  OAI2BB2XL U1871 ( .B0(n1141), .B1(n240), .A0N(M2[7]), .A1N(n240), .Y(n717)
         );
  OAI2BB2XL U1872 ( .B0(n1143), .B1(n241), .A0N(M1[0]), .A1N(n241), .Y(n718)
         );
  OAI2BB2XL U1873 ( .B0(n1143), .B1(n242), .A0N(M1[1]), .A1N(n242), .Y(n719)
         );
  OAI2BB2XL U1874 ( .B0(n1143), .B1(n243), .A0N(M1[2]), .A1N(n243), .Y(n720)
         );
  OAI2BB2XL U1875 ( .B0(n1143), .B1(n244), .A0N(M1[3]), .A1N(n244), .Y(n721)
         );
  OAI2BB2XL U1876 ( .B0(n1143), .B1(n245), .A0N(M1[4]), .A1N(n245), .Y(n722)
         );
  OAI2BB2XL U1877 ( .B0(n1143), .B1(n246), .A0N(M1[5]), .A1N(n246), .Y(n723)
         );
  OAI2BB2XL U1878 ( .B0(n1143), .B1(n247), .A0N(M1[6]), .A1N(n247), .Y(n724)
         );
  OAI2BB2XL U1879 ( .B0(n1143), .B1(n248), .A0N(M1[7]), .A1N(n248), .Y(n725)
         );
  CLKINVX1 U1880 ( .A(gray_data[1]), .Y(n1241) );
  CLKINVX1 U1881 ( .A(gray_data[0]), .Y(n1242) );
  CLKINVX1 U1882 ( .A(gray_valid), .Y(n1240) );
  CLKINVX1 U1883 ( .A(\SET[1][0] ), .Y(n1307) );
  CLKINVX1 U1884 ( .A(\SET[1][6] ), .Y(n1337) );
  CLKINVX1 U1885 ( .A(\SET[1][5] ), .Y(n1332) );
  CLKINVX1 U1886 ( .A(\SET[1][3] ), .Y(n1322) );
  CLKINVX1 U1887 ( .A(\SET[2][0] ), .Y(n1308) );
  NAND2BX1 U1888 ( .AN(n1136), .B(n629), .Y(n911) );
  NAND3X1 U1889 ( .A(n193), .B(n1151), .C(CNT_valid), .Y(n629) );
  OAI222XL U1890 ( .A0(n604), .A1(n1149), .B0(n594), .B1(n1253), .C0(n601), 
        .C1(num[0]), .Y(n603) );
  AO22X1 U1891 ( .A0(n627), .A1(amount[6]), .B0(N953), .B1(n628), .Y(n910) );
  AO22X1 U1892 ( .A0(n627), .A1(amount[5]), .B0(N952), .B1(n628), .Y(n904) );
  AO22X1 U1893 ( .A0(amount[4]), .A1(n627), .B0(N951), .B1(n628), .Y(n905) );
  AO22X1 U1894 ( .A0(amount[3]), .A1(n627), .B0(N950), .B1(n628), .Y(n906) );
  AO22X1 U1895 ( .A0(n627), .A1(amount[2]), .B0(N949), .B1(n628), .Y(n907) );
  AO22X1 U1896 ( .A0(amount[1]), .A1(n627), .B0(N948), .B1(n628), .Y(n908) );
  AO22X1 U1897 ( .A0(amount[0]), .A1(n627), .B0(N947), .B1(n628), .Y(n909) );
  CLKBUFX3 U1898 ( .A(N822), .Y(n1125) );
  OAI211X1 U1899 ( .A0(n1266), .A1(n84), .B0(n657), .C0(n658), .Y(N822) );
  AOI222XL U1900 ( .A0(\SET[3][6] ), .A1(n1267), .B0(\SET[5][6] ), .B1(n1268), 
        .C0(\SET[4][6] ), .C1(n1264), .Y(n658) );
  CLKINVX1 U1901 ( .A(\SET[1][7] ), .Y(n1341) );
  CLKINVX1 U1902 ( .A(\SET[2][7] ), .Y(n1342) );
  CLKINVX1 U1903 ( .A(\SET[2][6] ), .Y(n1338) );
  NAND2X1 U1904 ( .A(times[1]), .B(times[0]), .Y(n638) );
  NAND2X1 U1905 ( .A(times[2]), .B(n1254), .Y(n197) );
  CLKINVX1 U1906 ( .A(n638), .Y(n1254) );
  AOI222XL U1907 ( .A0(n1248), .A1(\SET_flag[3][1] ), .B0(n1250), .B1(
        \SET_flag[5][1] ), .C0(n1064), .C1(\SET_flag[4][1] ), .Y(n494) );
  AOI222XL U1908 ( .A0(n1248), .A1(\SET_flag[3][3] ), .B0(n1250), .B1(
        \SET_flag[5][3] ), .C0(n1064), .C1(\SET_flag[4][3] ), .Y(n484) );
  AOI222XL U1909 ( .A0(n1248), .A1(\SET_flag[3][4] ), .B0(n1250), .B1(
        \SET_flag[5][4] ), .C0(n1064), .C1(\SET_flag[4][4] ), .Y(n479) );
  AOI222XL U1910 ( .A0(n1248), .A1(\SET_flag[3][5] ), .B0(n1250), .B1(
        \SET_flag[5][5] ), .C0(n1064), .C1(\SET_flag[4][5] ), .Y(n469) );
  MXI2X1 U1911 ( .A(n1081), .B(n1096), .S0(n1121), .Y(N1784) );
  MXI3X1 U1912 ( .A(\SET[1][0] ), .B(\SET[3][0] ), .C(\SET[5][0] ), .S0(n1119), 
        .S1(n1116), .Y(n1096) );
  MXI3X1 U1913 ( .A(n1307), .B(n1080), .C(n1081), .S0(n1116), .S1(n1121), .Y(
        N1785) );
  MXI2X1 U1914 ( .A(\SET[3][0] ), .B(\SET[5][0] ), .S0(n1120), .Y(n1080) );
  NAND2X1 U1915 ( .A(n1137), .B(n81), .Y(n559) );
  NAND2X1 U1916 ( .A(\bitpos[5][2] ), .B(n258), .Y(n260) );
  NAND2X1 U1917 ( .A(\bitpos[4][2] ), .B(n273), .Y(n275) );
  NAND2X1 U1918 ( .A(\bitpos[3][2] ), .B(n288), .Y(n290) );
  NAND2X1 U1919 ( .A(\bitpos[2][2] ), .B(n303), .Y(n305) );
  NAND2X1 U1920 ( .A(\bitpos[1][2] ), .B(n318), .Y(n320) );
  NAND2X1 U1921 ( .A(\bitpos[0][2] ), .B(n333), .Y(n335) );
  MXI3X1 U1922 ( .A(\SET[0][0] ), .B(\SET[2][0] ), .C(\SET[4][0] ), .S0(n1119), 
        .S1(n1117), .Y(n1081) );
  MXI3X1 U1923 ( .A(\SET[0][1] ), .B(\SET[2][1] ), .C(\SET[4][1] ), .S0(n1119), 
        .S1(n1117), .Y(n1083) );
  MXI3X1 U1924 ( .A(\SET[0][2] ), .B(\SET[2][2] ), .C(\SET[4][2] ), .S0(n1119), 
        .S1(n1137), .Y(n1085) );
  MXI3X1 U1925 ( .A(\SET[0][3] ), .B(\SET[2][3] ), .C(\SET[4][3] ), .S0(n1119), 
        .S1(n1137), .Y(n1087) );
  MXI3X1 U1926 ( .A(\SET[0][4] ), .B(\SET[2][4] ), .C(\SET[4][4] ), .S0(n1119), 
        .S1(n1117), .Y(n1089) );
  MXI2X1 U1927 ( .A(\SET[3][1] ), .B(\SET[5][1] ), .S0(n1120), .Y(n1082) );
  MXI2X1 U1928 ( .A(\SET[3][2] ), .B(\SET[5][2] ), .S0(n1119), .Y(n1084) );
  MXI2X1 U1929 ( .A(\SET[3][3] ), .B(\SET[5][3] ), .S0(n1120), .Y(n1086) );
  MXI3X1 U1930 ( .A(\SET[1][1] ), .B(\SET[3][1] ), .C(\SET[5][1] ), .S0(n1118), 
        .S1(n1116), .Y(n1097) );
  INVX3 U1931 ( .A(endpoint[2]), .Y(n1138) );
  MXI2X1 U1932 ( .A(n1085), .B(n1098), .S0(n1121), .Y(N1782) );
  MXI3X1 U1933 ( .A(n1317), .B(n1084), .C(n1085), .S0(n1116), .S1(n1121), .Y(
        N1787) );
  MXI3X1 U1934 ( .A(\SET[1][2] ), .B(\SET[3][2] ), .C(\SET[5][2] ), .S0(n1118), 
        .S1(n1116), .Y(n1098) );
  MXI2X1 U1935 ( .A(n1087), .B(n1099), .S0(n1121), .Y(N1781) );
  MXI3X1 U1936 ( .A(n1322), .B(n1086), .C(n1087), .S0(n1116), .S1(n1121), .Y(
        N1788) );
  MXI3X1 U1937 ( .A(\SET[1][3] ), .B(\SET[3][3] ), .C(\SET[5][3] ), .S0(n1118), 
        .S1(n1116), .Y(n1099) );
  MXI2X1 U1938 ( .A(n1089), .B(n1100), .S0(n1132), .Y(N1780) );
  MXI3X1 U1939 ( .A(n1327), .B(n1088), .C(n1089), .S0(n1116), .S1(n1121), .Y(
        N1789) );
  MXI3X1 U1940 ( .A(\SET[1][4] ), .B(\SET[3][4] ), .C(\SET[5][4] ), .S0(n1118), 
        .S1(n1116), .Y(n1100) );
  MXI2X1 U1941 ( .A(n1091), .B(n1101), .S0(n1132), .Y(N1779) );
  MXI3X1 U1942 ( .A(n1332), .B(n1090), .C(n1091), .S0(n1116), .S1(n1121), .Y(
        N1790) );
  MXI3X1 U1943 ( .A(\SET[1][5] ), .B(\SET[3][5] ), .C(\SET[5][5] ), .S0(n1118), 
        .S1(n1117), .Y(n1101) );
  MXI2X1 U1944 ( .A(n1093), .B(n1102), .S0(n1132), .Y(N1778) );
  MXI3X1 U1945 ( .A(n1337), .B(n1092), .C(n1093), .S0(n1117), .S1(n1121), .Y(
        N1791) );
  MXI3X1 U1946 ( .A(\SET[1][6] ), .B(\SET[3][6] ), .C(\SET[5][6] ), .S0(n1118), 
        .S1(endpoint[2]), .Y(n1102) );
  CLKBUFX3 U1947 ( .A(n249), .Y(n1127) );
  OAI22XL U1948 ( .A0(n371), .A1(n1133), .B0(n1132), .B1(n372), .Y(n249) );
  AOI222XL U1949 ( .A0(\SET_flag[4][5] ), .A1(n1060), .B0(\SET_flag[0][5] ), 
        .B1(n1063), .C0(\SET_flag[2][5] ), .C1(n1261), .Y(n371) );
  AOI222XL U1950 ( .A0(\SET_flag[5][5] ), .A1(n1060), .B0(\SET_flag[1][5] ), 
        .B1(n1063), .C0(\SET_flag[3][5] ), .C1(n1261), .Y(n372) );
  CLKBUFX3 U1951 ( .A(n264), .Y(n1128) );
  OAI22XL U1952 ( .A0(n365), .A1(n1133), .B0(n1132), .B1(n366), .Y(n264) );
  AOI222XL U1953 ( .A0(\SET_flag[4][4] ), .A1(n1060), .B0(\SET_flag[0][4] ), 
        .B1(n1063), .C0(\SET_flag[2][4] ), .C1(n1261), .Y(n365) );
  AOI222XL U1954 ( .A0(\SET_flag[5][4] ), .A1(n1060), .B0(\SET_flag[1][4] ), 
        .B1(n1063), .C0(\SET_flag[3][4] ), .C1(n1261), .Y(n366) );
  CLKBUFX3 U1955 ( .A(n279), .Y(n1129) );
  OAI22XL U1956 ( .A0(n359), .A1(n1133), .B0(n1132), .B1(n360), .Y(n279) );
  AOI222XL U1957 ( .A0(\SET_flag[4][3] ), .A1(n1060), .B0(\SET_flag[0][3] ), 
        .B1(n1063), .C0(\SET_flag[2][3] ), .C1(n1261), .Y(n359) );
  AOI222XL U1958 ( .A0(\SET_flag[5][3] ), .A1(n1060), .B0(\SET_flag[1][3] ), 
        .B1(n1063), .C0(\SET_flag[3][3] ), .C1(n1261), .Y(n360) );
  CLKBUFX3 U1959 ( .A(n294), .Y(n1130) );
  OAI22XL U1960 ( .A0(n353), .A1(n1133), .B0(n1132), .B1(n354), .Y(n294) );
  AOI222XL U1961 ( .A0(\SET_flag[4][2] ), .A1(n1060), .B0(\SET_flag[0][2] ), 
        .B1(n1063), .C0(\SET_flag[2][2] ), .C1(n1261), .Y(n353) );
  AOI222XL U1962 ( .A0(\SET_flag[5][2] ), .A1(n1060), .B0(\SET_flag[1][2] ), 
        .B1(n1063), .C0(\SET_flag[3][2] ), .C1(n1261), .Y(n354) );
  CLKBUFX3 U1963 ( .A(n309), .Y(n1131) );
  OAI22XL U1964 ( .A0(n345), .A1(n1133), .B0(n1132), .B1(n346), .Y(n309) );
  AOI222XL U1965 ( .A0(\SET_flag[4][1] ), .A1(n1060), .B0(\SET_flag[0][1] ), 
        .B1(n1063), .C0(\SET_flag[2][1] ), .C1(n1261), .Y(n345) );
  AOI222XL U1966 ( .A0(\SET_flag[5][1] ), .A1(n1060), .B0(\SET_flag[1][1] ), 
        .B1(n1063), .C0(\SET_flag[3][1] ), .C1(n1261), .Y(n346) );
  CLKBUFX3 U1967 ( .A(n324), .Y(n1126) );
  OAI22XL U1968 ( .A0(n375), .A1(n1133), .B0(n1132), .B1(n376), .Y(n324) );
  AOI222XL U1969 ( .A0(\SET_flag[4][0] ), .A1(n1060), .B0(\SET_flag[0][0] ), 
        .B1(n1063), .C0(\SET_flag[2][0] ), .C1(n1261), .Y(n375) );
  AOI222XL U1970 ( .A0(\SET_flag[5][0] ), .A1(n1060), .B0(\SET_flag[1][0] ), 
        .B1(n1063), .C0(\SET_flag[3][0] ), .C1(n1261), .Y(n376) );
  CLKBUFX3 U1971 ( .A(endpoint[0]), .Y(n1132) );
  AOI222XL U1972 ( .A0(n1248), .A1(\SET_flag[3][2] ), .B0(n1250), .B1(
        \SET_flag[5][2] ), .C0(n1064), .C1(\SET_flag[4][2] ), .Y(n489) );
  OAI211X1 U1973 ( .A0(n1295), .A1(n1266), .B0(n495), .C0(n496), .Y(n399) );
  AOI222XL U1974 ( .A0(n1267), .A1(\SET_flag[3][1] ), .B0(n1268), .B1(
        \SET_flag[5][1] ), .C0(n1264), .C1(\SET_flag[4][1] ), .Y(n496) );
  OAI211X1 U1975 ( .A0(n1289), .A1(n1266), .B0(n490), .C0(n491), .Y(n395) );
  AOI222XL U1976 ( .A0(n1267), .A1(\SET_flag[3][2] ), .B0(n1268), .B1(
        \SET_flag[5][2] ), .C0(n1264), .C1(\SET_flag[4][2] ), .Y(n491) );
  OAI211X1 U1977 ( .A0(n1283), .A1(n1266), .B0(n485), .C0(n486), .Y(n391) );
  AOI222XL U1978 ( .A0(n1267), .A1(\SET_flag[3][3] ), .B0(n1268), .B1(
        \SET_flag[5][3] ), .C0(n1264), .C1(\SET_flag[4][3] ), .Y(n486) );
  OAI211X1 U1979 ( .A0(n1277), .A1(n1266), .B0(n480), .C0(n481), .Y(n387) );
  AOI222XL U1980 ( .A0(n1267), .A1(\SET_flag[3][4] ), .B0(n1268), .B1(
        \SET_flag[5][4] ), .C0(n1264), .C1(\SET_flag[4][4] ), .Y(n481) );
  OAI211X1 U1981 ( .A0(n1271), .A1(n1266), .B0(n472), .C0(n473), .Y(n383) );
  AOI222XL U1982 ( .A0(n1267), .A1(\SET_flag[3][5] ), .B0(n1268), .B1(
        \SET_flag[5][5] ), .C0(n1264), .C1(\SET_flag[4][5] ), .Y(n473) );
  OAI211X1 U1983 ( .A0(n1301), .A1(n1266), .B0(n498), .C0(n499), .Y(n404) );
  AOI222XL U1984 ( .A0(n1267), .A1(\SET_flag[3][0] ), .B0(n1268), .B1(
        \SET_flag[5][0] ), .C0(n1264), .C1(\SET_flag[4][0] ), .Y(n499) );
  MXI2X1 U1985 ( .A(n1069), .B(n1104), .S0(endpoint[0]), .Y(N840) );
  MXI3X1 U1986 ( .A(\SET_flag[1][0] ), .B(\SET_flag[3][0] ), .C(
        \SET_flag[5][0] ), .S0(n1118), .S1(n1117), .Y(n1104) );
  MXI2X1 U1987 ( .A(n1071), .B(n1105), .S0(endpoint[0]), .Y(N839) );
  MXI3X1 U1988 ( .A(\SET_flag[1][1] ), .B(\SET_flag[3][1] ), .C(
        \SET_flag[5][1] ), .S0(n1118), .S1(n1117), .Y(n1105) );
  MXI2X1 U1989 ( .A(n1073), .B(n1106), .S0(endpoint[0]), .Y(N838) );
  MXI3X1 U1990 ( .A(\SET_flag[1][2] ), .B(\SET_flag[3][2] ), .C(
        \SET_flag[5][2] ), .S0(n1118), .S1(n1137), .Y(n1106) );
  MXI2X1 U1991 ( .A(n1075), .B(n1107), .S0(endpoint[0]), .Y(N837) );
  MXI3X1 U1992 ( .A(\SET_flag[1][3] ), .B(\SET_flag[3][3] ), .C(
        \SET_flag[5][3] ), .S0(n1118), .S1(endpoint[2]), .Y(n1107) );
  MXI2X1 U1993 ( .A(n1077), .B(n1108), .S0(endpoint[0]), .Y(N836) );
  MXI3X1 U1994 ( .A(\SET_flag[1][4] ), .B(\SET_flag[3][4] ), .C(
        \SET_flag[5][4] ), .S0(n1118), .S1(n1116), .Y(n1108) );
  MXI2X1 U1995 ( .A(n1079), .B(n1109), .S0(n1132), .Y(N835) );
  MXI3X1 U1996 ( .A(\SET_flag[1][5] ), .B(\SET_flag[3][5] ), .C(
        \SET_flag[5][5] ), .S0(n1119), .S1(n1116), .Y(n1109) );
  NOR3X1 U1997 ( .A(state[1]), .B(state[2]), .C(n69), .Y(n630) );
  NOR3X1 U1998 ( .A(state[1]), .B(state[2]), .C(state[0]), .Y(n198) );
  MXI3X1 U1999 ( .A(\SET[0][5] ), .B(\SET[2][5] ), .C(\SET[4][5] ), .S0(n1119), 
        .S1(n1117), .Y(n1091) );
  MXI3X1 U2000 ( .A(\SET_flag[0][0] ), .B(\SET_flag[2][0] ), .C(
        \SET_flag[4][0] ), .S0(n1119), .S1(n1117), .Y(n1069) );
  MXI3X1 U2001 ( .A(\SET[0][6] ), .B(\SET[2][6] ), .C(\SET[4][6] ), .S0(n1119), 
        .S1(endpoint[2]), .Y(n1093) );
  MXI3X1 U2002 ( .A(\SET_flag[0][1] ), .B(\SET_flag[2][1] ), .C(
        \SET_flag[4][1] ), .S0(n1119), .S1(n1117), .Y(n1071) );
  MXI3X1 U2003 ( .A(\SET_flag[0][2] ), .B(\SET_flag[2][2] ), .C(
        \SET_flag[4][2] ), .S0(n1119), .S1(n1117), .Y(n1073) );
  MXI3X1 U2004 ( .A(\SET_flag[0][3] ), .B(\SET_flag[2][3] ), .C(
        \SET_flag[4][3] ), .S0(n1119), .S1(n1117), .Y(n1075) );
  MXI3X1 U2005 ( .A(\SET_flag[0][4] ), .B(\SET_flag[2][4] ), .C(
        \SET_flag[4][4] ), .S0(n1119), .S1(n1117), .Y(n1077) );
  MXI3X1 U2006 ( .A(\SET_flag[0][5] ), .B(\SET_flag[2][5] ), .C(
        \SET_flag[4][5] ), .S0(n1119), .S1(n1117), .Y(n1079) );
  MXI3X1 U2007 ( .A(\SET[0][7] ), .B(\SET[2][7] ), .C(\SET[4][7] ), .S0(n1119), 
        .S1(endpoint[2]), .Y(n1095) );
  MXI3X1 U2008 ( .A(n1111), .B(n1070), .C(n1071), .S0(n1116), .S1(n1121), .Y(
        N1868) );
  MXI2X1 U2009 ( .A(\SET_flag[3][1] ), .B(\SET_flag[5][1] ), .S0(n1120), .Y(
        n1070) );
  MXI3X1 U2010 ( .A(n1112), .B(n1072), .C(n1073), .S0(n1116), .S1(n1121), .Y(
        N1869) );
  MXI2X1 U2011 ( .A(\SET_flag[3][2] ), .B(\SET_flag[5][2] ), .S0(n1120), .Y(
        n1072) );
  MXI3X1 U2012 ( .A(n1113), .B(n1074), .C(n1075), .S0(n1116), .S1(n1121), .Y(
        N1870) );
  MXI2X1 U2013 ( .A(\SET_flag[3][3] ), .B(\SET_flag[5][3] ), .S0(n1120), .Y(
        n1074) );
  MXI3X1 U2014 ( .A(n1114), .B(n1076), .C(n1077), .S0(n1116), .S1(n1121), .Y(
        N1871) );
  MXI2X1 U2015 ( .A(\SET_flag[3][4] ), .B(\SET_flag[5][4] ), .S0(n1120), .Y(
        n1076) );
  MXI3X1 U2016 ( .A(n1115), .B(n1078), .C(n1079), .S0(n1116), .S1(n1121), .Y(
        N1872) );
  MXI2X1 U2017 ( .A(\SET_flag[3][5] ), .B(\SET_flag[5][5] ), .S0(n1120), .Y(
        n1078) );
  AOI222XL U2018 ( .A0(n1248), .A1(\SET_flag[3][0] ), .B0(n1250), .B1(
        \SET_flag[5][0] ), .C0(n1064), .C1(\SET_flag[4][0] ), .Y(n501) );
  NOR2X1 U2019 ( .A(N1867), .B(N840), .Y(n403) );
  MXI3X1 U2020 ( .A(n1110), .B(n1068), .C(n1069), .S0(n1116), .S1(n1121), .Y(
        N1867) );
  MXI2X1 U2021 ( .A(\SET_flag[3][0] ), .B(\SET_flag[5][0] ), .S0(n1120), .Y(
        n1068) );
  MXI2X1 U2022 ( .A(\SET[3][4] ), .B(\SET[5][4] ), .S0(n1119), .Y(n1088) );
  MXI2X1 U2023 ( .A(\SET[3][5] ), .B(\SET[5][5] ), .S0(n1120), .Y(n1090) );
  MXI2X1 U2024 ( .A(\SET[3][6] ), .B(\SET[5][6] ), .S0(n1120), .Y(n1092) );
  MXI2X1 U2025 ( .A(\SET[3][7] ), .B(\SET[5][7] ), .S0(n1120), .Y(n1094) );
  CLKINVX1 U2026 ( .A(\SET_flag[0][0] ), .Y(n1301) );
  CLKINVX1 U2027 ( .A(\SET_flag[0][1] ), .Y(n1295) );
  CLKINVX1 U2028 ( .A(\SET_flag[0][2] ), .Y(n1289) );
  CLKINVX1 U2029 ( .A(\SET_flag[0][3] ), .Y(n1283) );
  CLKINVX1 U2030 ( .A(\SET_flag[0][4] ), .Y(n1277) );
  CLKINVX1 U2031 ( .A(\SET_flag[0][5] ), .Y(n1271) );
  MXI3X1 U2032 ( .A(\SET[1][7] ), .B(\SET[3][7] ), .C(\SET[5][7] ), .S0(n1118), 
        .S1(endpoint[2]), .Y(n1103) );
  CLKINVX1 U2033 ( .A(\SET_flag[2][1] ), .Y(n1294) );
  CLKINVX1 U2034 ( .A(\SET_flag[2][2] ), .Y(n1288) );
  CLKINVX1 U2035 ( .A(\SET_flag[2][3] ), .Y(n1282) );
  CLKINVX1 U2036 ( .A(\SET_flag[2][4] ), .Y(n1276) );
  CLKINVX1 U2037 ( .A(\SET_flag[2][5] ), .Y(n1270) );
  OAI221XL U2038 ( .A0(n195), .A1(n196), .B0(n193), .B1(n197), .C0(n68), .Y(
        nextstate[0]) );
  OR4X1 U2039 ( .A(amount[0]), .B(amount[1]), .C(amount[3]), .D(amount[4]), 
        .Y(n195) );
  NAND4X1 U2040 ( .A(amount[6]), .B(amount[5]), .C(amount[2]), .D(n198), .Y(
        n196) );
  NAND3X1 U2041 ( .A(n81), .B(n1138), .C(n1132), .Y(n191) );
  NOR3X1 U2042 ( .A(n1138), .B(n1132), .C(n81), .Y(n466) );
  CLKINVX1 U2043 ( .A(\bitpos[0][0] ), .Y(n1303) );
  CLKINVX1 U2044 ( .A(\bitpos[5][0] ), .Y(n1273) );
  CLKINVX1 U2045 ( .A(\bitpos[4][0] ), .Y(n1279) );
  CLKINVX1 U2046 ( .A(\bitpos[3][0] ), .Y(n1285) );
  CLKINVX1 U2047 ( .A(\bitpos[2][0] ), .Y(n1291) );
  CLKINVX1 U2048 ( .A(\bitpos[1][0] ), .Y(n1297) );
  CLKINVX1 U2049 ( .A(\bitpos[0][1] ), .Y(n1304) );
  CLKINVX1 U2050 ( .A(\bitpos[5][1] ), .Y(n1274) );
  CLKINVX1 U2051 ( .A(\bitpos[4][1] ), .Y(n1280) );
  CLKINVX1 U2052 ( .A(\bitpos[3][1] ), .Y(n1286) );
  CLKINVX1 U2053 ( .A(\bitpos[2][1] ), .Y(n1292) );
  CLKINVX1 U2054 ( .A(\bitpos[1][1] ), .Y(n1298) );
  NAND2X1 U2055 ( .A(\bitpos[5][1] ), .B(n1273), .Y(n256) );
  NAND2X1 U2056 ( .A(\bitpos[4][1] ), .B(n1279), .Y(n271) );
  NAND2X1 U2057 ( .A(\bitpos[3][1] ), .B(n1285), .Y(n286) );
  NAND2X1 U2058 ( .A(\bitpos[2][1] ), .B(n1291), .Y(n301) );
  NAND2X1 U2059 ( .A(\bitpos[1][1] ), .B(n1297), .Y(n316) );
  NAND2X1 U2060 ( .A(\bitpos[0][1] ), .B(n1303), .Y(n331) );
  NAND2X1 U2061 ( .A(\bitpos[5][0] ), .B(n1274), .Y(n254) );
  NAND2X1 U2062 ( .A(\bitpos[4][0] ), .B(n1280), .Y(n269) );
  NAND2X1 U2063 ( .A(\bitpos[3][0] ), .B(n1286), .Y(n284) );
  NAND2X1 U2064 ( .A(\bitpos[2][0] ), .B(n1292), .Y(n299) );
  NAND2X1 U2065 ( .A(\bitpos[1][0] ), .B(n1298), .Y(n314) );
  NAND2X1 U2066 ( .A(\bitpos[0][0] ), .B(n1304), .Y(n329) );
  OAI21XL U2067 ( .A0(n191), .A1(n192), .B0(n68), .Y(nextstate[2]) );
  CLKINVX1 U2068 ( .A(times[0]), .Y(n1253) );
  NOR2X1 U2069 ( .A(times[1]), .B(times[0]), .Y(n637) );
  NAND3X1 U2070 ( .A(n193), .B(n1256), .C(n194), .Y(nextstate[1]) );
  NAND3X1 U2071 ( .A(n191), .B(n68), .C(state[0]), .Y(n194) );
  CLKINVX1 U2072 ( .A(\SET_flag[2][0] ), .Y(n1300) );
  CLKINVX1 U2073 ( .A(\bitpos[5][2] ), .Y(n1275) );
  CLKINVX1 U2074 ( .A(\bitpos[4][2] ), .Y(n1281) );
  CLKINVX1 U2075 ( .A(\bitpos[3][2] ), .Y(n1287) );
  CLKINVX1 U2076 ( .A(\bitpos[2][2] ), .Y(n1293) );
  CLKINVX1 U2077 ( .A(\bitpos[1][2] ), .Y(n1299) );
  CLKINVX1 U2078 ( .A(\bitpos[0][2] ), .Y(n1305) );
  CLKINVX1 U2079 ( .A(times[1]), .Y(n1262) );
  NAND2BX1 U2080 ( .AN(N810), .B(N824), .Y(n1168) );
  OAI222XL U2081 ( .A0(n1122), .A1(n1183), .B0(n1122), .B1(n1168), .C0(n1183), 
        .C1(n1168), .Y(n1169) );
  OAI222XL U2082 ( .A0(n1125), .A1(n1169), .B0(n1186), .B1(n1169), .C0(n1125), 
        .C1(n1186), .Y(n1180) );
  OAI22XL U2083 ( .A0(n1123), .A1(n1184), .B0(n1123), .B1(n1172), .Y(n1178) );
  NOR2BX1 U2084 ( .AN(N812), .B(N826), .Y(n1170) );
  OA22X1 U2085 ( .A0(n1170), .A1(n1123), .B0(n1170), .B1(n1184), .Y(n1174) );
  AOI21X1 U2086 ( .A0(N813), .A1(n1185), .B0(N814), .Y(n1171) );
  AOI2BB2X1 U2087 ( .B0(n1171), .B1(N828), .A0N(N813), .A1N(n1185), .Y(n1173)
         );
  OAI22XL U2088 ( .A0(n1175), .A1(n1183), .B0(n1122), .B1(n1175), .Y(n1176) );
  AO22X1 U2089 ( .A0(n1182), .A1(N807), .B0(n1180), .B1(n1179), .Y(n1181) );
  OAI21XL U2090 ( .A0(N807), .A1(n1182), .B0(n1181), .Y(N962) );
endmodule

